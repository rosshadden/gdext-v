module gd

pub enum CollisionObject3DDisableMode as i64 {
	disable_mode_remove = 0
	disable_mode_make_static = 1
	disable_mode_keep_active = 2
}

pub struct CollisionObject3D {
	Node3D
}

pub fn (s &CollisionObject3D) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s CollisionObject3D) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub interface ICollisionObject3DInputEvent {
mut:
	input_event_(camera Camera3D, event InputEvent, event_position Vector3, normal Vector3, shape_idx i64)
}

pub fn (s &CollisionObject3D) gd_input_event(camera Camera3D, event InputEvent, event_position Vector3, normal Vector3, shape_idx i64) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("_input_event")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2310605070)
	mut args := unsafe { [5]voidptr{} }
	args[0] = voidptr(&camera.ptr)
	args[1] = voidptr(&event.ptr)
	args[2] = unsafe{voidptr(&event_position)}
	args[3] = unsafe{voidptr(&normal)}
	args[4] = unsafe{voidptr(&shape_idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub interface ICollisionObject3DMouseEnter {
mut:
	mouse_enter_()
}

pub fn (s &CollisionObject3D) gd_mouse_enter() {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("_mouse_enter")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub interface ICollisionObject3DMouseExit {
mut:
	mouse_exit_()
}

pub fn (s &CollisionObject3D) gd_mouse_exit() {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("_mouse_exit")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) set_collision_layer(layer i64) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_collision_layer")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&layer)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_collision_layer() i64 {
	mut result := i64(0)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_collision_layer")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) set_collision_mask(mask i64) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_collision_mask")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&mask)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_collision_mask() i64 {
	mut result := i64(0)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_collision_mask")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) set_collision_layer_value(layer_number i64, value bool) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_collision_layer_value")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 300928843)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&layer_number)}
	args[1] = unsafe{voidptr(&value)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_collision_layer_value(layer_number i64) bool {
	mut result := false
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_collision_layer_value")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1116898809)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&layer_number)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) set_collision_mask_value(layer_number i64, value bool) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_collision_mask_value")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 300928843)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&layer_number)}
	args[1] = unsafe{voidptr(&value)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_collision_mask_value(layer_number i64) bool {
	mut result := false
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_collision_mask_value")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1116898809)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&layer_number)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) set_collision_priority(priority f64) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_collision_priority")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&priority)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_collision_priority() f64 {
	mut result := f64(0)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_collision_priority")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) set_disable_mode(mode CollisionObject3DDisableMode) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_disable_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1623620376)
	mut args := unsafe { [1]voidptr{} }
	i64_mode := i64(mode)
	args[0] = unsafe{voidptr(&i64_mode)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_disable_mode() CollisionObject3DDisableMode {
	mut result := i64(CollisionObject3DDisableMode.disable_mode_remove)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_disable_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 410164780)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return unsafe{CollisionObject3DDisableMode(result)}
}

pub fn (s &CollisionObject3D) set_ray_pickable(ray_pickable bool) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_ray_pickable")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&ray_pickable)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) is_ray_pickable() bool {
	mut result := false
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("is_ray_pickable")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) set_capture_input_on_drag(enable bool) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("set_capture_input_on_drag")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&enable)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_capture_input_on_drag() bool {
	mut result := false
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_capture_input_on_drag")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) get_rid() RID {
	mut result := RID{}
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_rid")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2944877500)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) create_shape_owner(owner Object) i64 {
	mut result := i64(0)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("create_shape_owner")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3429307534)
	mut args := unsafe { [1]voidptr{} }
	args[0] = voidptr(&owner.ptr)
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) remove_shape_owner(owner_id i64) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("remove_shape_owner")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) get_shape_owners() PackedInt32Array {
	mut result := PackedInt32Array{}
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("get_shape_owners")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 969006518)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) shape_owner_set_transform(owner_id i64, transform Transform3D) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_set_transform")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3616898986)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	args[1] = unsafe{voidptr(&transform)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) shape_owner_get_transform(owner_id i64) Transform3D {
	mut result := Transform3D{}
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_get_transform")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1965739696)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) shape_owner_get_owner(owner_id i64) Object {
	mut result := Object{}
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_get_owner")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3332903315)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) shape_owner_set_disabled(owner_id i64, disabled bool) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_set_disabled")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 300928843)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	args[1] = unsafe{voidptr(&disabled)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) is_shape_owner_disabled(owner_id i64) bool {
	mut result := false
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("is_shape_owner_disabled")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1116898809)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) shape_owner_add_shape(owner_id i64, shape Shape3D) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_add_shape")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2566676345)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	args[1] = voidptr(&shape.ptr)
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) shape_owner_get_shape_count(owner_id i64) i64 {
	mut result := i64(0)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_get_shape_count")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 923996154)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) shape_owner_get_shape(owner_id i64, shape_id i64) Shape3D {
	mut result := Shape3D{}
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_get_shape")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 4015519174)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	args[1] = unsafe{voidptr(&shape_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) shape_owner_get_shape_index(owner_id i64, shape_id i64) i64 {
	mut result := i64(0)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_get_shape_index")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3175239445)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	args[1] = unsafe{voidptr(&shape_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &CollisionObject3D) shape_owner_remove_shape(owner_id i64, shape_id i64) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_remove_shape")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3937882851)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	args[1] = unsafe{voidptr(&shape_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) shape_owner_clear_shapes(owner_id i64) {
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_owner_clear_shapes")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&owner_id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &CollisionObject3D) shape_find_owner(shape_index i64) i64 {
	mut result := i64(0)
	classname := StringName.new("CollisionObject3D")
	fnname := StringName.new("shape_find_owner")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 923996154)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&shape_index)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
