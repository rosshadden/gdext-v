module gd

pub struct AudioStreamPlaybackInteractive {
	AudioStreamPlayback
}

pub fn (s &AudioStreamPlaybackInteractive) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s AudioStreamPlaybackInteractive) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &AudioStreamPlaybackInteractive) switch_to_clip_by_name(clip_name string) {
	classname := StringName.new("AudioStreamPlaybackInteractive")
	fnname := StringName.new("switch_to_clip_by_name")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3304788590)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := StringName.new(clip_name)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
}

pub fn (s &AudioStreamPlaybackInteractive) switch_to_clip(clip_index i64) {
	classname := StringName.new("AudioStreamPlaybackInteractive")
	fnname := StringName.new("switch_to_clip")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&clip_index)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &AudioStreamPlaybackInteractive) get_current_clip_index() i64 {
	mut result := i64(0)
	classname := StringName.new("AudioStreamPlaybackInteractive")
	fnname := StringName.new("get_current_clip_index")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
