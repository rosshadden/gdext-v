module gd

pub enum DirectionalLight3DShadowMode as i64 {
	shadow_orthogonal = 0
	shadow_parallel_2_splits = 1
	shadow_parallel_4_splits = 2
}

pub enum DirectionalLight3DSkyMode as i64 {
	sky_mode_light_and_sky = 0
	sky_mode_light_only = 1
	sky_mode_sky_only = 2
}

pub struct DirectionalLight3D {
	Light3D
}

pub fn (s &DirectionalLight3D) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s DirectionalLight3D) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &DirectionalLight3D) set_shadow_mode(mode DirectionalLight3DShadowMode) {
	classname := StringName.new("DirectionalLight3D")
	fnname := StringName.new("set_shadow_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1261211726)
	mut args := unsafe { [1]voidptr{} }
	i64_mode := i64(mode)
	args[0] = unsafe{voidptr(&i64_mode)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &DirectionalLight3D) get_shadow_mode() DirectionalLight3DShadowMode {
	mut result := i64(DirectionalLight3DShadowMode.shadow_orthogonal)
	classname := StringName.new("DirectionalLight3D")
	fnname := StringName.new("get_shadow_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2765228544)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return unsafe{DirectionalLight3DShadowMode(result)}
}

pub fn (s &DirectionalLight3D) set_blend_splits(enabled bool) {
	classname := StringName.new("DirectionalLight3D")
	fnname := StringName.new("set_blend_splits")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&enabled)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &DirectionalLight3D) is_blend_splits_enabled() bool {
	mut result := false
	classname := StringName.new("DirectionalLight3D")
	fnname := StringName.new("is_blend_splits_enabled")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &DirectionalLight3D) set_sky_mode(mode DirectionalLight3DSkyMode) {
	classname := StringName.new("DirectionalLight3D")
	fnname := StringName.new("set_sky_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2691194817)
	mut args := unsafe { [1]voidptr{} }
	i64_mode := i64(mode)
	args[0] = unsafe{voidptr(&i64_mode)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &DirectionalLight3D) get_sky_mode() DirectionalLight3DSkyMode {
	mut result := i64(DirectionalLight3DSkyMode.sky_mode_light_and_sky)
	classname := StringName.new("DirectionalLight3D")
	fnname := StringName.new("get_sky_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3819982774)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return unsafe{DirectionalLight3DSkyMode(result)}
}
