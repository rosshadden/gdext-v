module gd

pub struct VisualShaderNodeParticleMultiplyByAxisAngle {
	VisualShaderNode
}

pub fn (s &VisualShaderNodeParticleMultiplyByAxisAngle) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s VisualShaderNodeParticleMultiplyByAxisAngle) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &VisualShaderNodeParticleMultiplyByAxisAngle) set_degrees_mode(enabled bool) {
	classname := StringName.new("VisualShaderNodeParticleMultiplyByAxisAngle")
	fnname := StringName.new("set_degrees_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&enabled)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &VisualShaderNodeParticleMultiplyByAxisAngle) is_degrees_mode() bool {
	mut result := false
	classname := StringName.new("VisualShaderNodeParticleMultiplyByAxisAngle")
	fnname := StringName.new("is_degrees_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
