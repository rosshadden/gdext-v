module gd

pub struct WorldBoundaryShape2D {
	Shape2D
}

pub fn (s &WorldBoundaryShape2D) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s WorldBoundaryShape2D) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &WorldBoundaryShape2D) set_normal(normal Vector2) {
	classname := StringName.new("WorldBoundaryShape2D")
	fnname := StringName.new("set_normal")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 743155724)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&normal)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &WorldBoundaryShape2D) get_normal() Vector2 {
	mut result := Vector2{}
	classname := StringName.new("WorldBoundaryShape2D")
	fnname := StringName.new("get_normal")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &WorldBoundaryShape2D) set_distance(distance f64) {
	classname := StringName.new("WorldBoundaryShape2D")
	fnname := StringName.new("set_distance")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&distance)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &WorldBoundaryShape2D) get_distance() f64 {
	mut result := f64(0)
	classname := StringName.new("WorldBoundaryShape2D")
	fnname := StringName.new("get_distance")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
