module gd

fn astar2d_gd_estimate_cost[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAStar2DEstimateCost(unsafe{&T(voidptr(inst))})
	from_id := unsafe{&i64(args[0])}
	end_id := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.estimate_cost_(from_id, end_id)
}

fn astar2d_gd_compute_cost[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAStar2DComputeCost(unsafe{&T(voidptr(inst))})
	from_id := unsafe{&i64(args[0])}
	to_id := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.compute_cost_(from_id, to_id)
}

fn astar3d_gd_estimate_cost[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAStar3DEstimateCost(unsafe{&T(voidptr(inst))})
	from_id := unsafe{&i64(args[0])}
	end_id := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.estimate_cost_(from_id, end_id)
}

fn astar3d_gd_compute_cost[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAStar3DComputeCost(unsafe{&T(voidptr(inst))})
	from_id := unsafe{&i64(args[0])}
	to_id := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.compute_cost_(from_id, to_id)
}

fn astargrid2d_gd_estimate_cost[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAStarGrid2DEstimateCost(unsafe{&T(voidptr(inst))})
	from_id := unsafe{&Vector2i(args[0])}
	end_id := unsafe{&Vector2i(args[1])}
	*(&f64(ret)) := v_inst.estimate_cost_(from_id, end_id)
}

fn astargrid2d_gd_compute_cost[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAStarGrid2DComputeCost(unsafe{&T(voidptr(inst))})
	from_id := unsafe{&Vector2i(args[0])}
	to_id := unsafe{&Vector2i(args[1])}
	*(&f64(ret)) := v_inst.compute_cost_(from_id, to_id)
}

fn animationmixer_gd_post_process_key_value[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationMixerPostProcessKeyValue(unsafe{&T(voidptr(inst))})
	animation := unsafe{&Animation(args[0])}
	track := unsafe{&i64(args[1])}
	value := unsafe{&Variant(args[2])}
	object_id := unsafe{&i64(args[3])}
	object_sub_idx := unsafe{&i64(args[4])}
	*(&Variant(ret)) := v_inst.post_process_key_value_(animation, track, value, object_id, object_sub_idx)
}

fn animationnode_gd_get_child_nodes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeGetChildNodes(unsafe{&T(voidptr(inst))})
	*(&Dictionary(ret)) := v_inst.get_child_nodes_()
}

fn animationnode_gd_get_parameter_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeGetParameterList(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_parameter_list_()
}

fn animationnode_gd_get_child_by_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeGetChildByName(unsafe{&T(voidptr(inst))})
	name := unsafe{&StringName(args[0])}
	*(&AnimationNode(ret)) := v_inst.get_child_by_name_(name)
}

fn animationnode_gd_get_parameter_default_value[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeGetParameterDefaultValue(unsafe{&T(voidptr(inst))})
	parameter := unsafe{&StringName(args[0])}
	*(&Variant(ret)) := v_inst.get_parameter_default_value_(parameter)
}

fn animationnode_gd_is_parameter_read_only[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeIsParameterReadOnly(unsafe{&T(voidptr(inst))})
	parameter := unsafe{&StringName(args[0])}
	*(&bool(ret)) := v_inst.is_parameter_read_only_(parameter)
}

fn animationnode_gd_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeProcess(unsafe{&T(voidptr(inst))})
	time := unsafe{&f64(args[0])}
	seek := unsafe{&bool(args[1])}
	is_external_seeking := unsafe{&bool(args[2])}
	test_only := unsafe{&bool(args[3])}
	*(&f64(ret)) := v_inst.process_(time, seek, is_external_seeking, test_only)
}

fn animationnode_gd_get_caption[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeGetCaption(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_caption_()
}

fn animationnode_gd_has_filter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeHasFilter(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_filter_()
}

fn animationnodeextension_gd_process_animation_node[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAnimationNodeExtensionProcessAnimationNode(unsafe{&T(voidptr(inst))})
	playback_info := unsafe{&PackedFloat64Array(args[0])}
	test_only := unsafe{&bool(args[1])}
	*(&PackedFloat32Array(ret)) := v_inst.process_animation_node_(playback_info, test_only)
}

fn audioeffect_gd_instantiate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioEffectInstantiate(unsafe{&T(voidptr(inst))})
	*(&AudioEffectInstance(ret)) := v_inst.instantiate_()
}

fn audioeffectinstance_gd_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioEffectInstanceProcess(unsafe{&T(voidptr(inst))})
	src_buffer := unsafe{&voidptr(args[0])}
	dst_buffer := unsafe{&&AudioFrame(args[1])}
	frame_count := unsafe{&i64(args[2])}
	v_inst.process_(src_buffer, dst_buffer, frame_count)
}

fn audioeffectinstance_gd_process_silence[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioEffectInstanceProcessSilence(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.process_silence_()
}

fn audiostream_gd_instantiate_playback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamInstantiatePlayback(unsafe{&T(voidptr(inst))})
	*(&AudioStreamPlayback(ret)) := v_inst.instantiate_playback_()
}

fn audiostream_gd_get_stream_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamGetStreamName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_stream_name_()
}

fn audiostream_gd_get_length[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamGetLength(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_length_()
}

fn audiostream_gd_is_monophonic[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamIsMonophonic(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_monophonic_()
}

fn audiostream_gd_get_bpm[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamGetBpm(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_bpm_()
}

fn audiostream_gd_get_beat_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamGetBeatCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_beat_count_()
}

fn audiostream_gd_get_parameter_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamGetParameterList(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_parameter_list_()
}

fn audiostream_gd_has_loop[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamHasLoop(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_loop_()
}

fn audiostream_gd_get_bar_beats[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamGetBarBeats(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_bar_beats_()
}

fn audiostreamplayback_gd_start[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackStart(unsafe{&T(voidptr(inst))})
	from_pos := unsafe{&f64(args[0])}
	v_inst.start_(from_pos)
}

fn audiostreamplayback_gd_stop[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackStop(unsafe{&T(voidptr(inst))})
	v_inst.stop_()
}

fn audiostreamplayback_gd_is_playing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackIsPlaying(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_playing_()
}

fn audiostreamplayback_gd_get_loop_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackGetLoopCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_loop_count_()
}

fn audiostreamplayback_gd_get_playback_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackGetPlaybackPosition(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_playback_position_()
}

fn audiostreamplayback_gd_seek[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackSeek(unsafe{&T(voidptr(inst))})
	position := unsafe{&f64(args[0])}
	v_inst.seek_(position)
}

fn audiostreamplayback_gd_mix[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackMix(unsafe{&T(voidptr(inst))})
	buffer := unsafe{&&AudioFrame(args[0])}
	rate_scale := unsafe{&f64(args[1])}
	frames := unsafe{&i64(args[2])}
	*(&i64(ret)) := v_inst.mix_(buffer, rate_scale, frames)
}

fn audiostreamplayback_gd_tag_used_streams[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackTagUsedStreams(unsafe{&T(voidptr(inst))})
	v_inst.tag_used_streams_()
}

fn audiostreamplayback_gd_set_parameter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackSetParameter(unsafe{&T(voidptr(inst))})
	name := unsafe{&StringName(args[0])}
	value := unsafe{&Variant(args[1])}
	v_inst.set_parameter_(name, value)
}

fn audiostreamplayback_gd_get_parameter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackGetParameter(unsafe{&T(voidptr(inst))})
	name := unsafe{&StringName(args[0])}
	*(&Variant(ret)) := v_inst.get_parameter_(name)
}

fn audiostreamplaybackresampled_gd_mix_resampled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackResampledMixResampled(unsafe{&T(voidptr(inst))})
	dst_buffer := unsafe{&&AudioFrame(args[0])}
	frame_count := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.mix_resampled_(dst_buffer, frame_count)
}

fn audiostreamplaybackresampled_gd_get_stream_sampling_rate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IAudioStreamPlaybackResampledGetStreamSamplingRate(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_stream_sampling_rate_()
}

fn basebutton_gd_pressed[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IBaseButtonPressed(unsafe{&T(voidptr(inst))})
	v_inst.pressed_()
}

fn basebutton_gd_toggled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IBaseButtonToggled(unsafe{&T(voidptr(inst))})
	toggled_on := unsafe{&bool(args[0])}
	v_inst.toggled_(toggled_on)
}

fn camerafeed_gd_activate_feed[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICameraFeedActivateFeed(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.activate_feed_()
}

fn camerafeed_gd_deactivate_feed[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICameraFeedDeactivateFeed(unsafe{&T(voidptr(inst))})
	v_inst.deactivate_feed_()
}

fn canvasitem_gd_draw[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICanvasItemDraw(unsafe{&T(voidptr(inst))})
	v_inst.draw_()
}

fn codeedit_gd_confirm_code_completion[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICodeEditConfirmCodeCompletion(unsafe{&T(voidptr(inst))})
	replace := unsafe{&bool(args[0])}
	v_inst.confirm_code_completion_(replace)
}

fn codeedit_gd_request_code_completion[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICodeEditRequestCodeCompletion(unsafe{&T(voidptr(inst))})
	force := unsafe{&bool(args[0])}
	v_inst.request_code_completion_(force)
}

fn codeedit_gd_filter_code_completion_candidates[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICodeEditFilterCodeCompletionCandidates(unsafe{&T(voidptr(inst))})
	candidates := unsafe{&Array(args[0])}
	*(&Array(ret)) := v_inst.filter_code_completion_candidates_(candidates)
}

fn collisionobject2d_gd_input_event[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject2DInputEvent(unsafe{&T(voidptr(inst))})
	viewport := unsafe{&Viewport(args[0])}
	event := unsafe{&InputEvent(args[1])}
	shape_idx := unsafe{&i64(args[2])}
	v_inst.input_event_(viewport, event, shape_idx)
}

fn collisionobject2d_gd_mouse_enter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject2DMouseEnter(unsafe{&T(voidptr(inst))})
	v_inst.mouse_enter_()
}

fn collisionobject2d_gd_mouse_exit[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject2DMouseExit(unsafe{&T(voidptr(inst))})
	v_inst.mouse_exit_()
}

fn collisionobject2d_gd_mouse_shape_enter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject2DMouseShapeEnter(unsafe{&T(voidptr(inst))})
	shape_idx := unsafe{&i64(args[0])}
	v_inst.mouse_shape_enter_(shape_idx)
}

fn collisionobject2d_gd_mouse_shape_exit[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject2DMouseShapeExit(unsafe{&T(voidptr(inst))})
	shape_idx := unsafe{&i64(args[0])}
	v_inst.mouse_shape_exit_(shape_idx)
}

fn collisionobject3d_gd_input_event[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject3DInputEvent(unsafe{&T(voidptr(inst))})
	camera := unsafe{&Camera3D(args[0])}
	event := unsafe{&InputEvent(args[1])}
	event_position := unsafe{&Vector3(args[2])}
	normal := unsafe{&Vector3(args[3])}
	shape_idx := unsafe{&i64(args[4])}
	v_inst.input_event_(camera, event, event_position, normal, shape_idx)
}

fn collisionobject3d_gd_mouse_enter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject3DMouseEnter(unsafe{&T(voidptr(inst))})
	v_inst.mouse_enter_()
}

fn collisionobject3d_gd_mouse_exit[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICollisionObject3DMouseExit(unsafe{&T(voidptr(inst))})
	v_inst.mouse_exit_()
}

fn compositoreffect_gd_render_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ICompositorEffectRenderCallback(unsafe{&T(voidptr(inst))})
	effect_callback_type := unsafe{&i64(args[0])}
	render_data := unsafe{&RenderData(args[1])}
	v_inst.render_callback_(effect_callback_type, render_data)
}

fn container_gd_get_allowed_size_flags_horizontal[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IContainerGetAllowedSizeFlagsHorizontal(unsafe{&T(voidptr(inst))})
	*(&PackedInt32Array(ret)) := v_inst.get_allowed_size_flags_horizontal_()
}

fn container_gd_get_allowed_size_flags_vertical[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IContainerGetAllowedSizeFlagsVertical(unsafe{&T(voidptr(inst))})
	*(&PackedInt32Array(ret)) := v_inst.get_allowed_size_flags_vertical_()
}

fn control_gd_has_point[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlHasPoint(unsafe{&T(voidptr(inst))})
	point := unsafe{&Vector2(args[0])}
	*(&bool(ret)) := v_inst.has_point_(point)
}

fn control_gd_structured_text_parser[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlStructuredTextParser(unsafe{&T(voidptr(inst))})
	gd_args := unsafe{&Array(args[0])}
	text := unsafe{&String(args[1])}
	*(&Array(ret)) := v_inst.structured_text_parser_(gd_args, text)
}

fn control_gd_get_minimum_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlGetMinimumSize(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_minimum_size_()
}

fn control_gd_get_tooltip[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlGetTooltip(unsafe{&T(voidptr(inst))})
	at_position := unsafe{&Vector2(args[0])}
	*(&String(ret)) := v_inst.get_tooltip_(at_position)
}

fn control_gd_get_drag_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlGetDragData(unsafe{&T(voidptr(inst))})
	at_position := unsafe{&Vector2(args[0])}
	*(&Variant(ret)) := v_inst.get_drag_data_(at_position)
}

fn control_gd_can_drop_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlCanDropData(unsafe{&T(voidptr(inst))})
	at_position := unsafe{&Vector2(args[0])}
	data := unsafe{&Variant(args[1])}
	*(&bool(ret)) := v_inst.can_drop_data_(at_position, data)
}

fn control_gd_drop_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlDropData(unsafe{&T(voidptr(inst))})
	at_position := unsafe{&Vector2(args[0])}
	data := unsafe{&Variant(args[1])}
	v_inst.drop_data_(at_position, data)
}

fn control_gd_make_custom_tooltip[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlMakeCustomTooltip(unsafe{&T(voidptr(inst))})
	for_text := unsafe{&String(args[0])}
	*(&Object(ret)) := v_inst.make_custom_tooltip_(for_text)
}

fn control_gd_accessibility_get_contextual_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlAccessibilityGetContextualInfo(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.accessibility_get_contextual_info_()
}

fn control_gd_gui_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IControlGuiInput(unsafe{&T(voidptr(inst))})
	event := unsafe{&InputEvent(args[0])}
	v_inst.gui_input_(event)
}

fn editorcontextmenuplugin_gd_popup_menu[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorContextMenuPluginPopupMenu(unsafe{&T(voidptr(inst))})
	paths := unsafe{&PackedStringArray(args[0])}
	v_inst.popup_menu_(paths)
}

fn editordebuggerplugin_gd_setup_session[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorDebuggerPluginSetupSession(unsafe{&T(voidptr(inst))})
	session_id := unsafe{&i64(args[0])}
	v_inst.setup_session_(session_id)
}

fn editordebuggerplugin_gd_has_capture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorDebuggerPluginHasCapture(unsafe{&T(voidptr(inst))})
	capture := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.has_capture_(capture)
}

fn editordebuggerplugin_gd_capture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorDebuggerPluginCapture(unsafe{&T(voidptr(inst))})
	message := unsafe{&String(args[0])}
	data := unsafe{&Array(args[1])}
	session_id := unsafe{&i64(args[2])}
	*(&bool(ret)) := v_inst.capture_(message, data, session_id)
}

fn editordebuggerplugin_gd_goto_script_line[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorDebuggerPluginGotoScriptLine(unsafe{&T(voidptr(inst))})
	script := unsafe{&Script(args[0])}
	line := unsafe{&i64(args[1])}
	v_inst.goto_script_line_(script, line)
}

fn editordebuggerplugin_gd_breakpoints_cleared_in_tree[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorDebuggerPluginBreakpointsClearedInTree(unsafe{&T(voidptr(inst))})
	v_inst.breakpoints_cleared_in_tree_()
}

fn editordebuggerplugin_gd_breakpoint_set_in_tree[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorDebuggerPluginBreakpointSetInTree(unsafe{&T(voidptr(inst))})
	script := unsafe{&Script(args[0])}
	line := unsafe{&i64(args[1])}
	enabled := unsafe{&bool(args[2])}
	v_inst.breakpoint_set_in_tree_(script, line, enabled)
}

fn editorexportplatformextension_gd_get_preset_features[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetPresetFeatures(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	*(&PackedStringArray(ret)) := v_inst.get_preset_features_(preset)
}

fn editorexportplatformextension_gd_is_executable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionIsExecutable(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.is_executable_(path)
}

fn editorexportplatformextension_gd_get_export_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetExportOptions(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_export_options_()
}

fn editorexportplatformextension_gd_should_update_export_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionShouldUpdateExportOptions(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.should_update_export_options_()
}

fn editorexportplatformextension_gd_get_export_option_visibility[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetExportOptionVisibility(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	option := unsafe{&String(args[1])}
	*(&bool(ret)) := v_inst.get_export_option_visibility_(preset, option)
}

fn editorexportplatformextension_gd_get_export_option_warning[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetExportOptionWarning(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	option := unsafe{&StringName(args[1])}
	*(&String(ret)) := v_inst.get_export_option_warning_(preset, option)
}

fn editorexportplatformextension_gd_get_os_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetOsName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_os_name_()
}

fn editorexportplatformextension_gd_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_name_()
}

fn editorexportplatformextension_gd_get_logo[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetLogo(unsafe{&T(voidptr(inst))})
	*(&Texture2D(ret)) := v_inst.get_logo_()
}

fn editorexportplatformextension_gd_poll_export[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionPollExport(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.poll_export_()
}

fn editorexportplatformextension_gd_get_options_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetOptionsCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_options_count_()
}

fn editorexportplatformextension_gd_get_options_tooltip[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetOptionsTooltip(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_options_tooltip_()
}

fn editorexportplatformextension_gd_get_option_icon[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetOptionIcon(unsafe{&T(voidptr(inst))})
	device := unsafe{&i64(args[0])}
	*(&ImageTexture(ret)) := v_inst.get_option_icon_(device)
}

fn editorexportplatformextension_gd_get_option_label[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetOptionLabel(unsafe{&T(voidptr(inst))})
	device := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.get_option_label_(device)
}

fn editorexportplatformextension_gd_get_option_tooltip[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetOptionTooltip(unsafe{&T(voidptr(inst))})
	device := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.get_option_tooltip_(device)
}

fn editorexportplatformextension_gd_get_device_architecture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetDeviceArchitecture(unsafe{&T(voidptr(inst))})
	device := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.get_device_architecture_(device)
}

fn editorexportplatformextension_gd_cleanup[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionCleanup(unsafe{&T(voidptr(inst))})
	v_inst.cleanup_()
}

fn editorexportplatformextension_gd_run[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionRun(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	device := unsafe{&i64(args[1])}
	debug_flags := unsafe{&EditorExportPlatformDebugFlags(args[2])}
	*(&GDError(ret)) := v_inst.run_(preset, device, debug_flags)
}

fn editorexportplatformextension_gd_get_run_icon[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetRunIcon(unsafe{&T(voidptr(inst))})
	*(&Texture2D(ret)) := v_inst.get_run_icon_()
}

fn editorexportplatformextension_gd_can_export[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionCanExport(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&bool(ret)) := v_inst.can_export_(preset, debug)
}

fn editorexportplatformextension_gd_has_valid_export_configuration[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionHasValidExportConfiguration(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&bool(ret)) := v_inst.has_valid_export_configuration_(preset, debug)
}

fn editorexportplatformextension_gd_has_valid_project_configuration[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionHasValidProjectConfiguration(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	*(&bool(ret)) := v_inst.has_valid_project_configuration_(preset)
}

fn editorexportplatformextension_gd_get_binary_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetBinaryExtensions(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	*(&PackedStringArray(ret)) := v_inst.get_binary_extensions_(preset)
}

fn editorexportplatformextension_gd_export_project[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionExportProject(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	debug := unsafe{&bool(args[1])}
	path := unsafe{&String(args[2])}
	flags := unsafe{&EditorExportPlatformDebugFlags(args[3])}
	*(&GDError(ret)) := v_inst.export_project_(preset, debug, path, flags)
}

fn editorexportplatformextension_gd_export_pack[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionExportPack(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	debug := unsafe{&bool(args[1])}
	path := unsafe{&String(args[2])}
	flags := unsafe{&EditorExportPlatformDebugFlags(args[3])}
	*(&GDError(ret)) := v_inst.export_pack_(preset, debug, path, flags)
}

fn editorexportplatformextension_gd_export_zip[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionExportZip(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	debug := unsafe{&bool(args[1])}
	path := unsafe{&String(args[2])}
	flags := unsafe{&EditorExportPlatformDebugFlags(args[3])}
	*(&GDError(ret)) := v_inst.export_zip_(preset, debug, path, flags)
}

fn editorexportplatformextension_gd_export_pack_patch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionExportPackPatch(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	debug := unsafe{&bool(args[1])}
	path := unsafe{&String(args[2])}
	patches := unsafe{&PackedStringArray(args[3])}
	flags := unsafe{&EditorExportPlatformDebugFlags(args[4])}
	*(&GDError(ret)) := v_inst.export_pack_patch_(preset, debug, path, patches, flags)
}

fn editorexportplatformextension_gd_export_zip_patch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionExportZipPatch(unsafe{&T(voidptr(inst))})
	preset := unsafe{&EditorExportPreset(args[0])}
	debug := unsafe{&bool(args[1])}
	path := unsafe{&String(args[2])}
	patches := unsafe{&PackedStringArray(args[3])}
	flags := unsafe{&EditorExportPlatformDebugFlags(args[4])}
	*(&GDError(ret)) := v_inst.export_zip_patch_(preset, debug, path, patches, flags)
}

fn editorexportplatformextension_gd_get_platform_features[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetPlatformFeatures(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_platform_features_()
}

fn editorexportplatformextension_gd_get_debug_protocol[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPlatformExtensionGetDebugProtocol(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_debug_protocol_()
}

fn editorexportplugin_gd_export_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginExportFile(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	gd_type := unsafe{&String(args[1])}
	features := unsafe{&PackedStringArray(args[2])}
	v_inst.export_file_(path, gd_type, features)
}

fn editorexportplugin_gd_export_begin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginExportBegin(unsafe{&T(voidptr(inst))})
	features := unsafe{&PackedStringArray(args[0])}
	is_debug := unsafe{&bool(args[1])}
	path := unsafe{&String(args[2])}
	flags := unsafe{&i64(args[3])}
	v_inst.export_begin_(features, is_debug, path, flags)
}

fn editorexportplugin_gd_export_end[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginExportEnd(unsafe{&T(voidptr(inst))})
	v_inst.export_end_()
}

fn editorexportplugin_gd_begin_customize_resources[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginBeginCustomizeResources(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	features := unsafe{&PackedStringArray(args[1])}
	*(&bool(ret)) := v_inst.begin_customize_resources_(platform, features)
}

fn editorexportplugin_gd_customize_resource[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginCustomizeResource(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	path := unsafe{&String(args[1])}
	*(&Resource(ret)) := v_inst.customize_resource_(resource, path)
}

fn editorexportplugin_gd_begin_customize_scenes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginBeginCustomizeScenes(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	features := unsafe{&PackedStringArray(args[1])}
	*(&bool(ret)) := v_inst.begin_customize_scenes_(platform, features)
}

fn editorexportplugin_gd_customize_scene[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginCustomizeScene(unsafe{&T(voidptr(inst))})
	scene := unsafe{&Node(args[0])}
	path := unsafe{&String(args[1])}
	*(&Node(ret)) := v_inst.customize_scene_(scene, path)
}

fn editorexportplugin_gd_get_customization_configuration_hash[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetCustomizationConfigurationHash(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_customization_configuration_hash_()
}

fn editorexportplugin_gd_end_customize_scenes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginEndCustomizeScenes(unsafe{&T(voidptr(inst))})
	v_inst.end_customize_scenes_()
}

fn editorexportplugin_gd_end_customize_resources[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginEndCustomizeResources(unsafe{&T(voidptr(inst))})
	v_inst.end_customize_resources_()
}

fn editorexportplugin_gd_get_export_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetExportOptions(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	*(&Array(ret)) := v_inst.get_export_options_(platform)
}

fn editorexportplugin_gd_get_export_options_overrides[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetExportOptionsOverrides(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	*(&Dictionary(ret)) := v_inst.get_export_options_overrides_(platform)
}

fn editorexportplugin_gd_should_update_export_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginShouldUpdateExportOptions(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	*(&bool(ret)) := v_inst.should_update_export_options_(platform)
}

fn editorexportplugin_gd_get_export_option_visibility[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetExportOptionVisibility(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	option := unsafe{&String(args[1])}
	*(&bool(ret)) := v_inst.get_export_option_visibility_(platform, option)
}

fn editorexportplugin_gd_get_export_option_warning[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetExportOptionWarning(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	option := unsafe{&String(args[1])}
	*(&String(ret)) := v_inst.get_export_option_warning_(platform, option)
}

fn editorexportplugin_gd_get_export_features[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetExportFeatures(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&PackedStringArray(ret)) := v_inst.get_export_features_(platform, debug)
}

fn editorexportplugin_gd_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_name_()
}

fn editorexportplugin_gd_supports_platform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginSupportsPlatform(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	*(&bool(ret)) := v_inst.supports_platform_(platform)
}

fn editorexportplugin_gd_get_android_dependencies[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetAndroidDependencies(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&PackedStringArray(ret)) := v_inst.get_android_dependencies_(platform, debug)
}

fn editorexportplugin_gd_get_android_dependencies_maven_repos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetAndroidDependenciesMavenRepos(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&PackedStringArray(ret)) := v_inst.get_android_dependencies_maven_repos_(platform, debug)
}

fn editorexportplugin_gd_get_android_libraries[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetAndroidLibraries(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&PackedStringArray(ret)) := v_inst.get_android_libraries_(platform, debug)
}

fn editorexportplugin_gd_get_android_manifest_activity_element_contents[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetAndroidManifestActivityElementContents(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&String(ret)) := v_inst.get_android_manifest_activity_element_contents_(platform, debug)
}

fn editorexportplugin_gd_get_android_manifest_application_element_contents[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetAndroidManifestApplicationElementContents(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&String(ret)) := v_inst.get_android_manifest_application_element_contents_(platform, debug)
}

fn editorexportplugin_gd_get_android_manifest_element_contents[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginGetAndroidManifestElementContents(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	debug := unsafe{&bool(args[1])}
	*(&String(ret)) := v_inst.get_android_manifest_element_contents_(platform, debug)
}

fn editorexportplugin_gd_update_android_prebuilt_manifest[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorExportPluginUpdateAndroidPrebuiltManifest(unsafe{&T(voidptr(inst))})
	platform := unsafe{&EditorExportPlatform(args[0])}
	manifest_data := unsafe{&PackedByteArray(args[1])}
	*(&PackedByteArray(ret)) := v_inst.update_android_prebuilt_manifest_(platform, manifest_data)
}

fn editorfilesystemimportformatsupportquery_gd_is_active[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorFileSystemImportFormatSupportQueryIsActive(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_active_()
}

fn editorfilesystemimportformatsupportquery_gd_get_file_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorFileSystemImportFormatSupportQueryGetFileExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_file_extensions_()
}

fn editorfilesystemimportformatsupportquery_gd_query[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorFileSystemImportFormatSupportQueryQuery(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.query_()
}

fn editorimportplugin_gd_get_importer_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetImporterName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_importer_name_()
}

fn editorimportplugin_gd_get_visible_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetVisibleName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_visible_name_()
}

fn editorimportplugin_gd_get_preset_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetPresetCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_preset_count_()
}

fn editorimportplugin_gd_get_preset_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetPresetName(unsafe{&T(voidptr(inst))})
	preset_index := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.get_preset_name_(preset_index)
}

fn editorimportplugin_gd_get_recognized_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetRecognizedExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_recognized_extensions_()
}

fn editorimportplugin_gd_get_import_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetImportOptions(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	preset_index := unsafe{&i64(args[1])}
	*(&Array(ret)) := v_inst.get_import_options_(path, preset_index)
}

fn editorimportplugin_gd_get_save_extension[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetSaveExtension(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_save_extension_()
}

fn editorimportplugin_gd_get_resource_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetResourceType(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_resource_type_()
}

fn editorimportplugin_gd_get_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetPriority(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_priority_()
}

fn editorimportplugin_gd_get_import_order[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetImportOrder(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_import_order_()
}

fn editorimportplugin_gd_get_format_version[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetFormatVersion(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_format_version_()
}

fn editorimportplugin_gd_get_option_visibility[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginGetOptionVisibility(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	option_name := unsafe{&StringName(args[1])}
	options := unsafe{&Dictionary(args[2])}
	*(&bool(ret)) := v_inst.get_option_visibility_(path, option_name, options)
}

fn editorimportplugin_gd_import[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginImport(unsafe{&T(voidptr(inst))})
	source_file := unsafe{&String(args[0])}
	save_path := unsafe{&String(args[1])}
	options := unsafe{&Dictionary(args[2])}
	platform_variants := unsafe{&Array(args[3])}
	gen_files := unsafe{&Array(args[4])}
	*(&GDError(ret)) := v_inst.gd_import_(source_file, save_path, options, platform_variants, gen_files)
}

fn editorimportplugin_gd_can_import_threaded[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorImportPluginCanImportThreaded(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_import_threaded_()
}

fn editorinspectorplugin_gd_can_handle[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorInspectorPluginCanHandle(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	*(&bool(ret)) := v_inst.can_handle_(object)
}

fn editorinspectorplugin_gd_parse_begin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorInspectorPluginParseBegin(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	v_inst.parse_begin_(object)
}

fn editorinspectorplugin_gd_parse_category[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorInspectorPluginParseCategory(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	category := unsafe{&String(args[1])}
	v_inst.parse_category_(object, category)
}

fn editorinspectorplugin_gd_parse_group[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorInspectorPluginParseGroup(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	group := unsafe{&String(args[1])}
	v_inst.parse_group_(object, group)
}

fn editorinspectorplugin_gd_parse_property[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorInspectorPluginParseProperty(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	gd_type := unsafe{&VariantType(args[1])}
	name := unsafe{&String(args[2])}
	hint_type := unsafe{&PropertyHint(args[3])}
	hint_string := unsafe{&String(args[4])}
	usage_flags := unsafe{&PropertyUsageFlags(args[5])}
	wide := unsafe{&bool(args[6])}
	*(&bool(ret)) := v_inst.parse_property_(object, gd_type, name, hint_type, hint_string, usage_flags, wide)
}

fn editorinspectorplugin_gd_parse_end[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorInspectorPluginParseEnd(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	v_inst.parse_end_(object)
}

fn editornode3dgizmo_gd_redraw[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoRedraw(unsafe{&T(voidptr(inst))})
	v_inst.redraw_()
}

fn editornode3dgizmo_gd_get_handle_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoGetHandleName(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	secondary := unsafe{&bool(args[1])}
	*(&String(ret)) := v_inst.get_handle_name_(id, secondary)
}

fn editornode3dgizmo_gd_is_handle_highlighted[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoIsHandleHighlighted(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	secondary := unsafe{&bool(args[1])}
	*(&bool(ret)) := v_inst.is_handle_highlighted_(id, secondary)
}

fn editornode3dgizmo_gd_get_handle_value[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoGetHandleValue(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	secondary := unsafe{&bool(args[1])}
	*(&Variant(ret)) := v_inst.get_handle_value_(id, secondary)
}

fn editornode3dgizmo_gd_begin_handle_action[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoBeginHandleAction(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	secondary := unsafe{&bool(args[1])}
	v_inst.begin_handle_action_(id, secondary)
}

fn editornode3dgizmo_gd_set_handle[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoSetHandle(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	secondary := unsafe{&bool(args[1])}
	camera := unsafe{&Camera3D(args[2])}
	point := unsafe{&Vector2(args[3])}
	v_inst.set_handle_(id, secondary, camera, point)
}

fn editornode3dgizmo_gd_commit_handle[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoCommitHandle(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	secondary := unsafe{&bool(args[1])}
	restore := unsafe{&Variant(args[2])}
	cancel := unsafe{&bool(args[3])}
	v_inst.commit_handle_(id, secondary, restore, cancel)
}

fn editornode3dgizmo_gd_subgizmos_intersect_ray[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoSubgizmosIntersectRay(unsafe{&T(voidptr(inst))})
	camera := unsafe{&Camera3D(args[0])}
	point := unsafe{&Vector2(args[1])}
	*(&i64(ret)) := v_inst.subgizmos_intersect_ray_(camera, point)
}

fn editornode3dgizmo_gd_subgizmos_intersect_frustum[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoSubgizmosIntersectFrustum(unsafe{&T(voidptr(inst))})
	camera := unsafe{&Camera3D(args[0])}
	frustum := unsafe{&Array(args[1])}
	*(&PackedInt32Array(ret)) := v_inst.subgizmos_intersect_frustum_(camera, frustum)
}

fn editornode3dgizmo_gd_set_subgizmo_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoSetSubgizmoTransform(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	transform := unsafe{&Transform3D(args[1])}
	v_inst.set_subgizmo_transform_(id, transform)
}

fn editornode3dgizmo_gd_get_subgizmo_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoGetSubgizmoTransform(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	*(&Transform3D(ret)) := v_inst.get_subgizmo_transform_(id)
}

fn editornode3dgizmo_gd_commit_subgizmos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoCommitSubgizmos(unsafe{&T(voidptr(inst))})
	ids := unsafe{&PackedInt32Array(args[0])}
	restores := unsafe{&Array(args[1])}
	cancel := unsafe{&bool(args[2])}
	v_inst.commit_subgizmos_(ids, restores, cancel)
}

fn editornode3dgizmoplugin_gd_has_gizmo[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginHasGizmo(unsafe{&T(voidptr(inst))})
	for_node_3d := unsafe{&Node3D(args[0])}
	*(&bool(ret)) := v_inst.has_gizmo_(for_node_3d)
}

fn editornode3dgizmoplugin_gd_create_gizmo[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginCreateGizmo(unsafe{&T(voidptr(inst))})
	for_node_3d := unsafe{&Node3D(args[0])}
	*(&EditorNode3DGizmo(ret)) := v_inst.create_gizmo_(for_node_3d)
}

fn editornode3dgizmoplugin_gd_get_gizmo_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginGetGizmoName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_gizmo_name_()
}

fn editornode3dgizmoplugin_gd_get_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginGetPriority(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_priority_()
}

fn editornode3dgizmoplugin_gd_can_be_hidden[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginCanBeHidden(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_be_hidden_()
}

fn editornode3dgizmoplugin_gd_is_selectable_when_hidden[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginIsSelectableWhenHidden(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_selectable_when_hidden_()
}

fn editornode3dgizmoplugin_gd_redraw[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginRedraw(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	v_inst.redraw_(gizmo)
}

fn editornode3dgizmoplugin_gd_get_handle_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginGetHandleName(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	handle_id := unsafe{&i64(args[1])}
	secondary := unsafe{&bool(args[2])}
	*(&String(ret)) := v_inst.get_handle_name_(gizmo, handle_id, secondary)
}

fn editornode3dgizmoplugin_gd_is_handle_highlighted[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginIsHandleHighlighted(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	handle_id := unsafe{&i64(args[1])}
	secondary := unsafe{&bool(args[2])}
	*(&bool(ret)) := v_inst.is_handle_highlighted_(gizmo, handle_id, secondary)
}

fn editornode3dgizmoplugin_gd_get_handle_value[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginGetHandleValue(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	handle_id := unsafe{&i64(args[1])}
	secondary := unsafe{&bool(args[2])}
	*(&Variant(ret)) := v_inst.get_handle_value_(gizmo, handle_id, secondary)
}

fn editornode3dgizmoplugin_gd_begin_handle_action[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginBeginHandleAction(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	handle_id := unsafe{&i64(args[1])}
	secondary := unsafe{&bool(args[2])}
	v_inst.begin_handle_action_(gizmo, handle_id, secondary)
}

fn editornode3dgizmoplugin_gd_set_handle[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginSetHandle(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	handle_id := unsafe{&i64(args[1])}
	secondary := unsafe{&bool(args[2])}
	camera := unsafe{&Camera3D(args[3])}
	screen_pos := unsafe{&Vector2(args[4])}
	v_inst.set_handle_(gizmo, handle_id, secondary, camera, screen_pos)
}

fn editornode3dgizmoplugin_gd_commit_handle[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginCommitHandle(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	handle_id := unsafe{&i64(args[1])}
	secondary := unsafe{&bool(args[2])}
	restore := unsafe{&Variant(args[3])}
	cancel := unsafe{&bool(args[4])}
	v_inst.commit_handle_(gizmo, handle_id, secondary, restore, cancel)
}

fn editornode3dgizmoplugin_gd_subgizmos_intersect_ray[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginSubgizmosIntersectRay(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	camera := unsafe{&Camera3D(args[1])}
	screen_pos := unsafe{&Vector2(args[2])}
	*(&i64(ret)) := v_inst.subgizmos_intersect_ray_(gizmo, camera, screen_pos)
}

fn editornode3dgizmoplugin_gd_subgizmos_intersect_frustum[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginSubgizmosIntersectFrustum(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	camera := unsafe{&Camera3D(args[1])}
	frustum_planes := unsafe{&Array(args[2])}
	*(&PackedInt32Array(ret)) := v_inst.subgizmos_intersect_frustum_(gizmo, camera, frustum_planes)
}

fn editornode3dgizmoplugin_gd_get_subgizmo_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginGetSubgizmoTransform(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	subgizmo_id := unsafe{&i64(args[1])}
	*(&Transform3D(ret)) := v_inst.get_subgizmo_transform_(gizmo, subgizmo_id)
}

fn editornode3dgizmoplugin_gd_set_subgizmo_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginSetSubgizmoTransform(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	subgizmo_id := unsafe{&i64(args[1])}
	transform := unsafe{&Transform3D(args[2])}
	v_inst.set_subgizmo_transform_(gizmo, subgizmo_id, transform)
}

fn editornode3dgizmoplugin_gd_commit_subgizmos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorNode3DGizmoPluginCommitSubgizmos(unsafe{&T(voidptr(inst))})
	gizmo := unsafe{&EditorNode3DGizmo(args[0])}
	ids := unsafe{&PackedInt32Array(args[1])}
	restores := unsafe{&Array(args[2])}
	cancel := unsafe{&bool(args[3])}
	v_inst.commit_subgizmos_(gizmo, ids, restores, cancel)
}

fn editorplugin_gd_forward_canvas_gui_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginForwardCanvasGuiInput(unsafe{&T(voidptr(inst))})
	event := unsafe{&InputEvent(args[0])}
	*(&bool(ret)) := v_inst.forward_canvas_gui_input_(event)
}

fn editorplugin_gd_forward_canvas_draw_over_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginForwardCanvasDrawOverViewport(unsafe{&T(voidptr(inst))})
	viewport_control := unsafe{&Control(args[0])}
	v_inst.forward_canvas_draw_over_viewport_(viewport_control)
}

fn editorplugin_gd_forward_canvas_force_draw_over_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginForwardCanvasForceDrawOverViewport(unsafe{&T(voidptr(inst))})
	viewport_control := unsafe{&Control(args[0])}
	v_inst.forward_canvas_force_draw_over_viewport_(viewport_control)
}

fn editorplugin_gd_forward_3d_gui_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginForward3dGuiInput(unsafe{&T(voidptr(inst))})
	viewport_camera := unsafe{&Camera3D(args[0])}
	event := unsafe{&InputEvent(args[1])}
	*(&i64(ret)) := v_inst.forward_3d_gui_input_(viewport_camera, event)
}

fn editorplugin_gd_forward_3d_draw_over_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginForward3dDrawOverViewport(unsafe{&T(voidptr(inst))})
	viewport_control := unsafe{&Control(args[0])}
	v_inst.forward_3d_draw_over_viewport_(viewport_control)
}

fn editorplugin_gd_forward_3d_force_draw_over_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginForward3dForceDrawOverViewport(unsafe{&T(voidptr(inst))})
	viewport_control := unsafe{&Control(args[0])}
	v_inst.forward_3d_force_draw_over_viewport_(viewport_control)
}

fn editorplugin_gd_get_plugin_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginGetPluginName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_plugin_name_()
}

fn editorplugin_gd_get_plugin_icon[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginGetPluginIcon(unsafe{&T(voidptr(inst))})
	*(&Texture2D(ret)) := v_inst.get_plugin_icon_()
}

fn editorplugin_gd_has_main_screen[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginHasMainScreen(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_main_screen_()
}

fn editorplugin_gd_make_visible[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginMakeVisible(unsafe{&T(voidptr(inst))})
	visible := unsafe{&bool(args[0])}
	v_inst.make_visible_(visible)
}

fn editorplugin_gd_edit[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginEdit(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	v_inst.edit_(object)
}

fn editorplugin_gd_handles[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginHandles(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	*(&bool(ret)) := v_inst.handles_(object)
}

fn editorplugin_gd_get_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginGetState(unsafe{&T(voidptr(inst))})
	*(&Dictionary(ret)) := v_inst.get_state_()
}

fn editorplugin_gd_set_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginSetState(unsafe{&T(voidptr(inst))})
	state := unsafe{&Dictionary(args[0])}
	v_inst.set_state_(state)
}

fn editorplugin_gd_clear[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginClear(unsafe{&T(voidptr(inst))})
	v_inst.clear_()
}

fn editorplugin_gd_get_unsaved_status[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginGetUnsavedStatus(unsafe{&T(voidptr(inst))})
	for_scene := unsafe{&String(args[0])}
	*(&String(ret)) := v_inst.get_unsaved_status_(for_scene)
}

fn editorplugin_gd_save_external_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginSaveExternalData(unsafe{&T(voidptr(inst))})
	v_inst.save_external_data_()
}

fn editorplugin_gd_apply_changes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginApplyChanges(unsafe{&T(voidptr(inst))})
	v_inst.apply_changes_()
}

fn editorplugin_gd_get_breakpoints[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginGetBreakpoints(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_breakpoints_()
}

fn editorplugin_gd_set_window_layout[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginSetWindowLayout(unsafe{&T(voidptr(inst))})
	configuration := unsafe{&ConfigFile(args[0])}
	v_inst.set_window_layout_(configuration)
}

fn editorplugin_gd_get_window_layout[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginGetWindowLayout(unsafe{&T(voidptr(inst))})
	configuration := unsafe{&ConfigFile(args[0])}
	v_inst.get_window_layout_(configuration)
}

fn editorplugin_gd_build[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginBuild(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.build_()
}

fn editorplugin_gd_enable_plugin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginEnablePlugin(unsafe{&T(voidptr(inst))})
	v_inst.enable_plugin_()
}

fn editorplugin_gd_disable_plugin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPluginDisablePlugin(unsafe{&T(voidptr(inst))})
	v_inst.disable_plugin_()
}

fn editorproperty_gd_update_property[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPropertyUpdateProperty(unsafe{&T(voidptr(inst))})
	v_inst.update_property_()
}

fn editorproperty_gd_set_read_only[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorPropertySetReadOnly(unsafe{&T(voidptr(inst))})
	read_only := unsafe{&bool(args[0])}
	v_inst.set_read_only_(read_only)
}

fn editorresourceconversionplugin_gd_converts_to[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourceConversionPluginConvertsTo(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.converts_to_()
}

fn editorresourceconversionplugin_gd_handles[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourceConversionPluginHandles(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	*(&bool(ret)) := v_inst.handles_(resource)
}

fn editorresourceconversionplugin_gd_convert[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourceConversionPluginConvert(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	*(&Resource(ret)) := v_inst.convert_(resource)
}

fn editorresourcepicker_gd_set_create_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourcePickerSetCreateOptions(unsafe{&T(voidptr(inst))})
	menu_node := unsafe{&Object(args[0])}
	v_inst.set_create_options_(menu_node)
}

fn editorresourcepicker_gd_handle_menu_selected[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourcePickerHandleMenuSelected(unsafe{&T(voidptr(inst))})
	id := unsafe{&i64(args[0])}
	*(&bool(ret)) := v_inst.handle_menu_selected_(id)
}

fn editorresourcepreviewgenerator_gd_handles[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourcePreviewGeneratorHandles(unsafe{&T(voidptr(inst))})
	gd_type := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.handles_(gd_type)
}

fn editorresourcepreviewgenerator_gd_generate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourcePreviewGeneratorGenerate(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	size := unsafe{&Vector2i(args[1])}
	metadata := unsafe{&Dictionary(args[2])}
	*(&Texture2D(ret)) := v_inst.generate_(resource, size, metadata)
}

fn editorresourcepreviewgenerator_gd_generate_from_path[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourcePreviewGeneratorGenerateFromPath(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	size := unsafe{&Vector2i(args[1])}
	metadata := unsafe{&Dictionary(args[2])}
	*(&Texture2D(ret)) := v_inst.generate_from_path_(path, size, metadata)
}

fn editorresourcepreviewgenerator_gd_generate_small_preview_automatically[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourcePreviewGeneratorGenerateSmallPreviewAutomatically(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.generate_small_preview_automatically_()
}

fn editorresourcepreviewgenerator_gd_can_generate_small_preview[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourcePreviewGeneratorCanGenerateSmallPreview(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_generate_small_preview_()
}

fn editorresourcetooltipplugin_gd_handles[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourceTooltipPluginHandles(unsafe{&T(voidptr(inst))})
	gd_type := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.handles_(gd_type)
}

fn editorresourcetooltipplugin_gd_make_tooltip_for_path[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorResourceTooltipPluginMakeTooltipForPath(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	metadata := unsafe{&Dictionary(args[1])}
	base := unsafe{&Control(args[2])}
	*(&Control(ret)) := v_inst.make_tooltip_for_path_(path, metadata, base)
}

fn editorsceneformatimporter_gd_get_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorSceneFormatImporterGetExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_extensions_()
}

fn editorsceneformatimporter_gd_import_scene[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorSceneFormatImporterImportScene(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	flags := unsafe{&i64(args[1])}
	options := unsafe{&Dictionary(args[2])}
	*(&Object(ret)) := v_inst.import_scene_(path, flags, options)
}

fn editorsceneformatimporter_gd_get_import_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorSceneFormatImporterGetImportOptions(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	v_inst.get_import_options_(path)
}

fn editorsceneformatimporter_gd_get_option_visibility[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorSceneFormatImporterGetOptionVisibility(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	for_animation := unsafe{&bool(args[1])}
	option := unsafe{&String(args[2])}
	*(&Variant(ret)) := v_inst.get_option_visibility_(path, for_animation, option)
}

fn editorscenepostimport_gd_post_import[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPostImport(unsafe{&T(voidptr(inst))})
	scene := unsafe{&Node(args[0])}
	*(&Object(ret)) := v_inst.post_import_(scene)
}

fn editorscenepostimportplugin_gd_get_internal_import_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginGetInternalImportOptions(unsafe{&T(voidptr(inst))})
	category := unsafe{&i64(args[0])}
	v_inst.get_internal_import_options_(category)
}

fn editorscenepostimportplugin_gd_get_internal_option_visibility[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginGetInternalOptionVisibility(unsafe{&T(voidptr(inst))})
	category := unsafe{&i64(args[0])}
	for_animation := unsafe{&bool(args[1])}
	option := unsafe{&String(args[2])}
	*(&Variant(ret)) := v_inst.get_internal_option_visibility_(category, for_animation, option)
}

fn editorscenepostimportplugin_gd_get_internal_option_update_view_required[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginGetInternalOptionUpdateViewRequired(unsafe{&T(voidptr(inst))})
	category := unsafe{&i64(args[0])}
	option := unsafe{&String(args[1])}
	*(&Variant(ret)) := v_inst.get_internal_option_update_view_required_(category, option)
}

fn editorscenepostimportplugin_gd_internal_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginInternalProcess(unsafe{&T(voidptr(inst))})
	category := unsafe{&i64(args[0])}
	base_node := unsafe{&Node(args[1])}
	node := unsafe{&Node(args[2])}
	resource := unsafe{&Resource(args[3])}
	v_inst.internal_process_(category, base_node, node, resource)
}

fn editorscenepostimportplugin_gd_get_import_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginGetImportOptions(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	v_inst.get_import_options_(path)
}

fn editorscenepostimportplugin_gd_get_option_visibility[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginGetOptionVisibility(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	for_animation := unsafe{&bool(args[1])}
	option := unsafe{&String(args[2])}
	*(&Variant(ret)) := v_inst.get_option_visibility_(path, for_animation, option)
}

fn editorscenepostimportplugin_gd_pre_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginPreProcess(unsafe{&T(voidptr(inst))})
	scene := unsafe{&Node(args[0])}
	v_inst.pre_process_(scene)
}

fn editorscenepostimportplugin_gd_post_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScenePostImportPluginPostProcess(unsafe{&T(voidptr(inst))})
	scene := unsafe{&Node(args[0])}
	v_inst.post_process_(scene)
}

fn editorscript_gd_run[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorScriptRun(unsafe{&T(voidptr(inst))})
	v_inst.run_()
}

fn editorsyntaxhighlighter_gd_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorSyntaxHighlighterGetName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_name_()
}

fn editorsyntaxhighlighter_gd_get_supported_languages[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorSyntaxHighlighterGetSupportedLanguages(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_supported_languages_()
}

fn editortranslationparserplugin_gd_parse_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorTranslationParserPluginParseFile(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&Array(ret)) := v_inst.parse_file_(path)
}

fn editortranslationparserplugin_gd_get_recognized_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorTranslationParserPluginGetRecognizedExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_recognized_extensions_()
}

fn editorvcsinterface_gd_initialize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceInitialize(unsafe{&T(voidptr(inst))})
	project_path := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.initialize_(project_path)
}

fn editorvcsinterface_gd_set_credentials[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceSetCredentials(unsafe{&T(voidptr(inst))})
	username := unsafe{&String(args[0])}
	password := unsafe{&String(args[1])}
	ssh_public_key_path := unsafe{&String(args[2])}
	ssh_private_key_path := unsafe{&String(args[3])}
	ssh_passphrase := unsafe{&String(args[4])}
	v_inst.set_credentials_(username, password, ssh_public_key_path, ssh_private_key_path, ssh_passphrase)
}

fn editorvcsinterface_gd_get_modified_files_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetModifiedFilesData(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_modified_files_data_()
}

fn editorvcsinterface_gd_stage_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceStageFile(unsafe{&T(voidptr(inst))})
	file_path := unsafe{&String(args[0])}
	v_inst.stage_file_(file_path)
}

fn editorvcsinterface_gd_unstage_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceUnstageFile(unsafe{&T(voidptr(inst))})
	file_path := unsafe{&String(args[0])}
	v_inst.unstage_file_(file_path)
}

fn editorvcsinterface_gd_discard_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceDiscardFile(unsafe{&T(voidptr(inst))})
	file_path := unsafe{&String(args[0])}
	v_inst.discard_file_(file_path)
}

fn editorvcsinterface_gd_commit[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceCommit(unsafe{&T(voidptr(inst))})
	msg := unsafe{&String(args[0])}
	v_inst.commit_(msg)
}

fn editorvcsinterface_gd_get_diff[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetDiff(unsafe{&T(voidptr(inst))})
	identifier := unsafe{&String(args[0])}
	area := unsafe{&i64(args[1])}
	*(&Array(ret)) := v_inst.get_diff_(identifier, area)
}

fn editorvcsinterface_gd_shut_down[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceShutDown(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.shut_down_()
}

fn editorvcsinterface_gd_get_vcs_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetVcsName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_vcs_name_()
}

fn editorvcsinterface_gd_get_previous_commits[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetPreviousCommits(unsafe{&T(voidptr(inst))})
	max_commits := unsafe{&i64(args[0])}
	*(&Array(ret)) := v_inst.get_previous_commits_(max_commits)
}

fn editorvcsinterface_gd_get_branch_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetBranchList(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_branch_list_()
}

fn editorvcsinterface_gd_get_remotes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetRemotes(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_remotes_()
}

fn editorvcsinterface_gd_create_branch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceCreateBranch(unsafe{&T(voidptr(inst))})
	branch_name := unsafe{&String(args[0])}
	v_inst.create_branch_(branch_name)
}

fn editorvcsinterface_gd_remove_branch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceRemoveBranch(unsafe{&T(voidptr(inst))})
	branch_name := unsafe{&String(args[0])}
	v_inst.remove_branch_(branch_name)
}

fn editorvcsinterface_gd_create_remote[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceCreateRemote(unsafe{&T(voidptr(inst))})
	remote_name := unsafe{&String(args[0])}
	remote_url := unsafe{&String(args[1])}
	v_inst.create_remote_(remote_name, remote_url)
}

fn editorvcsinterface_gd_remove_remote[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceRemoveRemote(unsafe{&T(voidptr(inst))})
	remote_name := unsafe{&String(args[0])}
	v_inst.remove_remote_(remote_name)
}

fn editorvcsinterface_gd_get_current_branch_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetCurrentBranchName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_current_branch_name_()
}

fn editorvcsinterface_gd_checkout_branch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceCheckoutBranch(unsafe{&T(voidptr(inst))})
	branch_name := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.checkout_branch_(branch_name)
}

fn editorvcsinterface_gd_pull[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfacePull(unsafe{&T(voidptr(inst))})
	remote := unsafe{&String(args[0])}
	v_inst.pull_(remote)
}

fn editorvcsinterface_gd_push[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfacePush(unsafe{&T(voidptr(inst))})
	remote := unsafe{&String(args[0])}
	force := unsafe{&bool(args[1])}
	v_inst.push_(remote, force)
}

fn editorvcsinterface_gd_fetch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceFetch(unsafe{&T(voidptr(inst))})
	remote := unsafe{&String(args[0])}
	v_inst.fetch_(remote)
}

fn editorvcsinterface_gd_get_line_diff[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEditorVCSInterfaceGetLineDiff(unsafe{&T(voidptr(inst))})
	file_path := unsafe{&String(args[0])}
	text := unsafe{&String(args[1])}
	*(&Array(ret)) := v_inst.get_line_diff_(file_path, text)
}

fn engineprofiler_gd_toggle[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEngineProfilerToggle(unsafe{&T(voidptr(inst))})
	enable := unsafe{&bool(args[0])}
	options := unsafe{&Array(args[1])}
	v_inst.toggle_(enable, options)
}

fn engineprofiler_gd_add_frame[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEngineProfilerAddFrame(unsafe{&T(voidptr(inst))})
	data := unsafe{&Array(args[0])}
	v_inst.add_frame_(data)
}

fn engineprofiler_gd_tick[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IEngineProfilerTick(unsafe{&T(voidptr(inst))})
	frame_time := unsafe{&f64(args[0])}
	process_time := unsafe{&f64(args[1])}
	physics_time := unsafe{&f64(args[2])}
	physics_frame_time := unsafe{&f64(args[3])}
	v_inst.tick_(frame_time, process_time, physics_time, physics_frame_time)
}

fn gltfdocumentextension_gd_import_preflight[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionImportPreflight(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	extensions := unsafe{&PackedStringArray(args[1])}
	*(&GDError(ret)) := v_inst.import_preflight_(state, extensions)
}

fn gltfdocumentextension_gd_get_supported_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionGetSupportedExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_supported_extensions_()
}

fn gltfdocumentextension_gd_parse_node_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionParseNodeExtensions(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	gltf_node := unsafe{&GLTFNode(args[1])}
	extensions := unsafe{&Dictionary(args[2])}
	*(&GDError(ret)) := v_inst.parse_node_extensions_(state, gltf_node, extensions)
}

fn gltfdocumentextension_gd_parse_image_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionParseImageData(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	image_data := unsafe{&PackedByteArray(args[1])}
	mime_type := unsafe{&String(args[2])}
	ret_image := unsafe{&Image(args[3])}
	*(&GDError(ret)) := v_inst.parse_image_data_(state, image_data, mime_type, ret_image)
}

fn gltfdocumentextension_gd_get_image_file_extension[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionGetImageFileExtension(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_image_file_extension_()
}

fn gltfdocumentextension_gd_parse_texture_json[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionParseTextureJson(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	texture_json := unsafe{&Dictionary(args[1])}
	ret_gltf_texture := unsafe{&GLTFTexture(args[2])}
	*(&GDError(ret)) := v_inst.parse_texture_json_(state, texture_json, ret_gltf_texture)
}

fn gltfdocumentextension_gd_import_object_model_property[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionImportObjectModelProperty(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	split_json_pointer := unsafe{&PackedStringArray(args[1])}
	partial_paths := unsafe{&Array(args[2])}
	*(&GLTFObjectModelProperty(ret)) := v_inst.import_object_model_property_(state, split_json_pointer, partial_paths)
}

fn gltfdocumentextension_gd_import_post_parse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionImportPostParse(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	*(&GDError(ret)) := v_inst.import_post_parse_(state)
}

fn gltfdocumentextension_gd_import_pre_generate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionImportPreGenerate(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	*(&GDError(ret)) := v_inst.import_pre_generate_(state)
}

fn gltfdocumentextension_gd_generate_scene_node[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionGenerateSceneNode(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	gltf_node := unsafe{&GLTFNode(args[1])}
	scene_parent := unsafe{&Node(args[2])}
	*(&Node3D(ret)) := v_inst.generate_scene_node_(state, gltf_node, scene_parent)
}

fn gltfdocumentextension_gd_import_node[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionImportNode(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	gltf_node := unsafe{&GLTFNode(args[1])}
	json := unsafe{&Dictionary(args[2])}
	node := unsafe{&Node(args[3])}
	*(&GDError(ret)) := v_inst.import_node_(state, gltf_node, json, node)
}

fn gltfdocumentextension_gd_import_post[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionImportPost(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	root := unsafe{&Node(args[1])}
	*(&GDError(ret)) := v_inst.import_post_(state, root)
}

fn gltfdocumentextension_gd_export_preflight[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionExportPreflight(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	root := unsafe{&Node(args[1])}
	*(&GDError(ret)) := v_inst.export_preflight_(state, root)
}

fn gltfdocumentextension_gd_convert_scene_node[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionConvertSceneNode(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	gltf_node := unsafe{&GLTFNode(args[1])}
	scene_node := unsafe{&Node(args[2])}
	v_inst.convert_scene_node_(state, gltf_node, scene_node)
}

fn gltfdocumentextension_gd_export_post_convert[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionExportPostConvert(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	root := unsafe{&Node(args[1])}
	*(&GDError(ret)) := v_inst.export_post_convert_(state, root)
}

fn gltfdocumentextension_gd_export_preserialize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionExportPreserialize(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	*(&GDError(ret)) := v_inst.export_preserialize_(state)
}

fn gltfdocumentextension_gd_export_object_model_property[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionExportObjectModelProperty(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	node_path := unsafe{&NodePath(args[1])}
	godot_node := unsafe{&Node(args[2])}
	gltf_node_index := unsafe{&i64(args[3])}
	target_object := unsafe{&Object(args[4])}
	target_depth := unsafe{&i64(args[5])}
	*(&GLTFObjectModelProperty(ret)) := v_inst.export_object_model_property_(state, node_path, godot_node, gltf_node_index, target_object, target_depth)
}

fn gltfdocumentextension_gd_get_saveable_image_formats[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionGetSaveableImageFormats(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_saveable_image_formats_()
}

fn gltfdocumentextension_gd_serialize_image_to_bytes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionSerializeImageToBytes(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	image := unsafe{&Image(args[1])}
	image_dict := unsafe{&Dictionary(args[2])}
	image_format := unsafe{&String(args[3])}
	lossy_quality := unsafe{&f64(args[4])}
	*(&PackedByteArray(ret)) := v_inst.serialize_image_to_bytes_(state, image, image_dict, image_format, lossy_quality)
}

fn gltfdocumentextension_gd_save_image_at_path[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionSaveImageAtPath(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	image := unsafe{&Image(args[1])}
	file_path := unsafe{&String(args[2])}
	image_format := unsafe{&String(args[3])}
	lossy_quality := unsafe{&f64(args[4])}
	*(&GDError(ret)) := v_inst.save_image_at_path_(state, image, file_path, image_format, lossy_quality)
}

fn gltfdocumentextension_gd_serialize_texture_json[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionSerializeTextureJson(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	texture_json := unsafe{&Dictionary(args[1])}
	gltf_texture := unsafe{&GLTFTexture(args[2])}
	image_format := unsafe{&String(args[3])}
	*(&GDError(ret)) := v_inst.serialize_texture_json_(state, texture_json, gltf_texture, image_format)
}

fn gltfdocumentextension_gd_export_node[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionExportNode(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	gltf_node := unsafe{&GLTFNode(args[1])}
	json := unsafe{&Dictionary(args[2])}
	node := unsafe{&Node(args[3])}
	*(&GDError(ret)) := v_inst.export_node_(state, gltf_node, json, node)
}

fn gltfdocumentextension_gd_export_post[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGLTFDocumentExtensionExportPost(unsafe{&T(voidptr(inst))})
	state := unsafe{&GLTFState(args[0])}
	*(&GDError(ret)) := v_inst.export_post_(state)
}

fn graphedit_gd_is_in_input_hotzone[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGraphEditIsInInputHotzone(unsafe{&T(voidptr(inst))})
	in_node := unsafe{&Object(args[0])}
	in_port := unsafe{&i64(args[1])}
	mouse_position := unsafe{&Vector2(args[2])}
	*(&bool(ret)) := v_inst.is_in_input_hotzone_(in_node, in_port, mouse_position)
}

fn graphedit_gd_is_in_output_hotzone[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGraphEditIsInOutputHotzone(unsafe{&T(voidptr(inst))})
	in_node := unsafe{&Object(args[0])}
	in_port := unsafe{&i64(args[1])}
	mouse_position := unsafe{&Vector2(args[2])}
	*(&bool(ret)) := v_inst.is_in_output_hotzone_(in_node, in_port, mouse_position)
}

fn graphedit_gd_get_connection_line[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGraphEditGetConnectionLine(unsafe{&T(voidptr(inst))})
	from_position := unsafe{&Vector2(args[0])}
	to_position := unsafe{&Vector2(args[1])}
	*(&PackedVector2Array(ret)) := v_inst.get_connection_line_(from_position, to_position)
}

fn graphedit_gd_is_node_hover_valid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGraphEditIsNodeHoverValid(unsafe{&T(voidptr(inst))})
	from_node := unsafe{&StringName(args[0])}
	from_port := unsafe{&i64(args[1])}
	to_node := unsafe{&StringName(args[2])}
	to_port := unsafe{&i64(args[3])}
	*(&bool(ret)) := v_inst.is_node_hover_valid_(from_node, from_port, to_node, to_port)
}

fn graphnode_gd_draw_port[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IGraphNodeDrawPort(unsafe{&T(voidptr(inst))})
	slot_index := unsafe{&i64(args[0])}
	position := unsafe{&Vector2i(args[1])}
	left := unsafe{&bool(args[2])}
	color := unsafe{&Color(args[3])}
	v_inst.draw_port_(slot_index, position, left, color)
}

fn imageformatloaderextension_gd_get_recognized_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IImageFormatLoaderExtensionGetRecognizedExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_recognized_extensions_()
}

fn imageformatloaderextension_gd_load_image[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IImageFormatLoaderExtensionLoadImage(unsafe{&T(voidptr(inst))})
	image := unsafe{&Image(args[0])}
	fileaccess := unsafe{&FileAccess(args[1])}
	flags := unsafe{&ImageFormatLoaderLoaderFlags(args[2])}
	scale := unsafe{&f64(args[3])}
	*(&GDError(ret)) := v_inst.load_image_(image, fileaccess, flags, scale)
}

fn mainloop_gd_initialize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMainLoopInitialize(unsafe{&T(voidptr(inst))})
	v_inst.initialize_()
}

fn mainloop_gd_physics_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMainLoopPhysicsProcess(unsafe{&T(voidptr(inst))})
	delta := unsafe{&f64(args[0])}
	*(&bool(ret)) := v_inst.physics_process_(delta)
}

fn mainloop_gd_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMainLoopProcess(unsafe{&T(voidptr(inst))})
	delta := unsafe{&f64(args[0])}
	*(&bool(ret)) := v_inst.process_(delta)
}

fn mainloop_gd_finalize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMainLoopFinalize(unsafe{&T(voidptr(inst))})
	v_inst.finalize_()
}

fn material_gd_get_shader_rid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMaterialGetShaderRid(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_shader_rid_()
}

fn material_gd_get_shader_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMaterialGetShaderMode(unsafe{&T(voidptr(inst))})
	*(&ShaderMode(ret)) := v_inst.get_shader_mode_()
}

fn material_gd_can_do_next_pass[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMaterialCanDoNextPass(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_do_next_pass_()
}

fn material_gd_can_use_render_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMaterialCanUseRenderPriority(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_use_render_priority_()
}

fn mesh_gd_get_surface_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshGetSurfaceCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_surface_count_()
}

fn mesh_gd_surface_get_array_len[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetArrayLen(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.surface_get_array_len_(index)
}

fn mesh_gd_surface_get_array_index_len[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetArrayIndexLen(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.surface_get_array_index_len_(index)
}

fn mesh_gd_surface_get_arrays[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetArrays(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&Array(ret)) := v_inst.surface_get_arrays_(index)
}

fn mesh_gd_surface_get_blend_shape_arrays[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetBlendShapeArrays(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&Array(ret)) := v_inst.surface_get_blend_shape_arrays_(index)
}

fn mesh_gd_surface_get_lods[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetLods(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&Dictionary(ret)) := v_inst.surface_get_lods_(index)
}

fn mesh_gd_surface_get_format[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetFormat(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.surface_get_format_(index)
}

fn mesh_gd_surface_get_primitive_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetPrimitiveType(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.surface_get_primitive_type_(index)
}

fn mesh_gd_surface_set_material[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceSetMaterial(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	material := unsafe{&Material(args[1])}
	v_inst.surface_set_material_(index, material)
}

fn mesh_gd_surface_get_material[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSurfaceGetMaterial(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&Material(ret)) := v_inst.surface_get_material_(index)
}

fn mesh_gd_get_blend_shape_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshGetBlendShapeCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_blend_shape_count_()
}

fn mesh_gd_get_blend_shape_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshGetBlendShapeName(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&StringName(ret)) := v_inst.get_blend_shape_name_(index)
}

fn mesh_gd_set_blend_shape_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshSetBlendShapeName(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	name := unsafe{&StringName(args[1])}
	v_inst.set_blend_shape_name_(index, name)
}

fn mesh_gd_get_aabb[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMeshGetAabb(unsafe{&T(voidptr(inst))})
	*(&AABB(ret)) := v_inst.get_aabb_()
}

fn moviewriter_gd_get_audio_mix_rate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMovieWriterGetAudioMixRate(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_audio_mix_rate_()
}

fn moviewriter_gd_get_audio_speaker_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMovieWriterGetAudioSpeakerMode(unsafe{&T(voidptr(inst))})
	*(&AudioServerSpeakerMode(ret)) := v_inst.get_audio_speaker_mode_()
}

fn moviewriter_gd_handles_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMovieWriterHandlesFile(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.handles_file_(path)
}

fn moviewriter_gd_write_begin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMovieWriterWriteBegin(unsafe{&T(voidptr(inst))})
	movie_size := unsafe{&Vector2i(args[0])}
	fps := unsafe{&i64(args[1])}
	base_path := unsafe{&String(args[2])}
	*(&GDError(ret)) := v_inst.write_begin_(movie_size, fps, base_path)
}

fn moviewriter_gd_write_frame[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMovieWriterWriteFrame(unsafe{&T(voidptr(inst))})
	frame_image := unsafe{&Image(args[0])}
	audio_frame_block := unsafe{&voidptr(args[1])}
	*(&GDError(ret)) := v_inst.write_frame_(frame_image, audio_frame_block)
}

fn moviewriter_gd_write_end[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMovieWriterWriteEnd(unsafe{&T(voidptr(inst))})
	v_inst.write_end_()
}

fn multiplayerapiextension_gd_poll[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionPoll(unsafe{&T(voidptr(inst))})
	*(&GDError(ret)) := v_inst.poll_()
}

fn multiplayerapiextension_gd_set_multiplayer_peer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionSetMultiplayerPeer(unsafe{&T(voidptr(inst))})
	multiplayer_peer := unsafe{&MultiplayerPeer(args[0])}
	v_inst.set_multiplayer_peer_(multiplayer_peer)
}

fn multiplayerapiextension_gd_get_multiplayer_peer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionGetMultiplayerPeer(unsafe{&T(voidptr(inst))})
	*(&MultiplayerPeer(ret)) := v_inst.get_multiplayer_peer_()
}

fn multiplayerapiextension_gd_get_unique_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionGetUniqueId(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_unique_id_()
}

fn multiplayerapiextension_gd_get_peer_ids[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionGetPeerIds(unsafe{&T(voidptr(inst))})
	*(&PackedInt32Array(ret)) := v_inst.get_peer_ids_()
}

fn multiplayerapiextension_gd_rpc[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionRpc(unsafe{&T(voidptr(inst))})
	peer := unsafe{&i64(args[0])}
	object := unsafe{&Object(args[1])}
	method := unsafe{&StringName(args[2])}
	gd_args := unsafe{&Array(args[3])}
	*(&GDError(ret)) := v_inst.rpc_(peer, object, method, gd_args)
}

fn multiplayerapiextension_gd_get_remote_sender_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionGetRemoteSenderId(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_remote_sender_id_()
}

fn multiplayerapiextension_gd_object_configuration_add[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionObjectConfigurationAdd(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	configuration := unsafe{&Variant(args[1])}
	*(&GDError(ret)) := v_inst.object_configuration_add_(object, configuration)
}

fn multiplayerapiextension_gd_object_configuration_remove[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerAPIExtensionObjectConfigurationRemove(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	configuration := unsafe{&Variant(args[1])}
	*(&GDError(ret)) := v_inst.object_configuration_remove_(object, configuration)
}

fn multiplayerpeerextension_gd_get_packet[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetPacket(unsafe{&T(voidptr(inst))})
	r_buffer := unsafe{&&&u8 (args[0])}
	r_buffer_size := unsafe{&&i32(args[1])}
	*(&GDError(ret)) := v_inst.get_packet_(r_buffer, r_buffer_size)
}

fn multiplayerpeerextension_gd_put_packet[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionPutPacket(unsafe{&T(voidptr(inst))})
	p_buffer := unsafe{&&u8(args[0])}
	p_buffer_size := unsafe{&i64(args[1])}
	*(&GDError(ret)) := v_inst.put_packet_(p_buffer, p_buffer_size)
}

fn multiplayerpeerextension_gd_get_available_packet_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetAvailablePacketCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_available_packet_count_()
}

fn multiplayerpeerextension_gd_get_max_packet_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetMaxPacketSize(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_max_packet_size_()
}

fn multiplayerpeerextension_gd_get_packet_script[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetPacketScript(unsafe{&T(voidptr(inst))})
	*(&PackedByteArray(ret)) := v_inst.get_packet_script_()
}

fn multiplayerpeerextension_gd_put_packet_script[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionPutPacketScript(unsafe{&T(voidptr(inst))})
	p_buffer := unsafe{&PackedByteArray(args[0])}
	*(&GDError(ret)) := v_inst.put_packet_script_(p_buffer)
}

fn multiplayerpeerextension_gd_get_packet_channel[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetPacketChannel(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_packet_channel_()
}

fn multiplayerpeerextension_gd_get_packet_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetPacketMode(unsafe{&T(voidptr(inst))})
	*(&MultiplayerPeerTransferMode(ret)) := v_inst.get_packet_mode_()
}

fn multiplayerpeerextension_gd_set_transfer_channel[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionSetTransferChannel(unsafe{&T(voidptr(inst))})
	p_channel := unsafe{&i64(args[0])}
	v_inst.set_transfer_channel_(p_channel)
}

fn multiplayerpeerextension_gd_get_transfer_channel[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetTransferChannel(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_transfer_channel_()
}

fn multiplayerpeerextension_gd_set_transfer_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionSetTransferMode(unsafe{&T(voidptr(inst))})
	p_mode := unsafe{&MultiplayerPeerTransferMode(args[0])}
	v_inst.set_transfer_mode_(p_mode)
}

fn multiplayerpeerextension_gd_get_transfer_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetTransferMode(unsafe{&T(voidptr(inst))})
	*(&MultiplayerPeerTransferMode(ret)) := v_inst.get_transfer_mode_()
}

fn multiplayerpeerextension_gd_set_target_peer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionSetTargetPeer(unsafe{&T(voidptr(inst))})
	p_peer := unsafe{&i64(args[0])}
	v_inst.set_target_peer_(p_peer)
}

fn multiplayerpeerextension_gd_get_packet_peer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetPacketPeer(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_packet_peer_()
}

fn multiplayerpeerextension_gd_is_server[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionIsServer(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_server_()
}

fn multiplayerpeerextension_gd_poll[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionPoll(unsafe{&T(voidptr(inst))})
	v_inst.poll_()
}

fn multiplayerpeerextension_gd_close[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionClose(unsafe{&T(voidptr(inst))})
	v_inst.close_()
}

fn multiplayerpeerextension_gd_disconnect_peer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionDisconnectPeer(unsafe{&T(voidptr(inst))})
	p_peer := unsafe{&i64(args[0])}
	p_force := unsafe{&bool(args[1])}
	v_inst.disconnect_peer_(p_peer, p_force)
}

fn multiplayerpeerextension_gd_get_unique_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetUniqueId(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_unique_id_()
}

fn multiplayerpeerextension_gd_set_refuse_new_connections[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionSetRefuseNewConnections(unsafe{&T(voidptr(inst))})
	p_enable := unsafe{&bool(args[0])}
	v_inst.set_refuse_new_connections_(p_enable)
}

fn multiplayerpeerextension_gd_is_refusing_new_connections[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionIsRefusingNewConnections(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_refusing_new_connections_()
}

fn multiplayerpeerextension_gd_is_server_relay_supported[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionIsServerRelaySupported(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_server_relay_supported_()
}

fn multiplayerpeerextension_gd_get_connection_status[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IMultiplayerPeerExtensionGetConnectionStatus(unsafe{&T(voidptr(inst))})
	*(&MultiplayerPeerConnectionStatus(ret)) := v_inst.get_connection_status_()
}

fn node_gd_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeProcess(unsafe{&T(voidptr(inst))})
	delta := unsafe{&f64(args[0])}
	v_inst.process_(delta)
}

fn node_gd_physics_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodePhysicsProcess(unsafe{&T(voidptr(inst))})
	delta := unsafe{&f64(args[0])}
	v_inst.physics_process_(delta)
}

fn node_gd_enter_tree[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeEnterTree(unsafe{&T(voidptr(inst))})
	v_inst.enter_tree_()
}

fn node_gd_exit_tree[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeExitTree(unsafe{&T(voidptr(inst))})
	v_inst.exit_tree_()
}

fn node_gd_ready[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeReady(unsafe{&T(voidptr(inst))})
	v_inst.ready_()
}

fn node_gd_get_configuration_warnings[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeGetConfigurationWarnings(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_configuration_warnings_()
}

fn node_gd_get_accessibility_configuration_warnings[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeGetAccessibilityConfigurationWarnings(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_accessibility_configuration_warnings_()
}

fn node_gd_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeInput(unsafe{&T(voidptr(inst))})
	event := unsafe{&InputEvent(args[0])}
	v_inst.input_(event)
}

fn node_gd_shortcut_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeShortcutInput(unsafe{&T(voidptr(inst))})
	event := unsafe{&InputEvent(args[0])}
	v_inst.shortcut_input_(event)
}

fn node_gd_unhandled_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeUnhandledInput(unsafe{&T(voidptr(inst))})
	event := unsafe{&InputEvent(args[0])}
	v_inst.unhandled_input_(event)
}

fn node_gd_unhandled_key_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeUnhandledKeyInput(unsafe{&T(voidptr(inst))})
	event := unsafe{&InputEvent(args[0])}
	v_inst.unhandled_key_input_(event)
}

fn node_gd_get_focused_accessibility_element[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeGetFocusedAccessibilityElement(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_focused_accessibility_element_()
}

fn node_gd_get_accessibility_container_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &INodeGetAccessibilityContainerName(unsafe{&T(voidptr(inst))})
	node := unsafe{&Node(args[0])}
	*(&String(ret)) := v_inst.get_accessibility_container_name_(node)
}

fn openxrbindingmodifier_gd_get_description[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRBindingModifierGetDescription(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_description_()
}

fn openxrbindingmodifier_gd_get_ip_modification[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRBindingModifierGetIpModification(unsafe{&T(voidptr(inst))})
	*(&PackedByteArray(ret)) := v_inst.get_ip_modification_()
}

fn openxrextensionwrapper_gd_get_requested_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperGetRequestedExtensions(unsafe{&T(voidptr(inst))})
	*(&Dictionary(ret)) := v_inst.get_requested_extensions_()
}

fn openxrextensionwrapper_gd_set_system_properties_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetSystemPropertiesAndGetNextPointer(unsafe{&T(voidptr(inst))})
	next_pointer := unsafe{&voidptr(args[0])}
	*(&i64(ret)) := v_inst.set_system_properties_and_get_next_pointer_(next_pointer)
}

fn openxrextensionwrapper_gd_set_instance_create_info_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetInstanceCreateInfoAndGetNextPointer(unsafe{&T(voidptr(inst))})
	next_pointer := unsafe{&voidptr(args[0])}
	*(&i64(ret)) := v_inst.set_instance_create_info_and_get_next_pointer_(next_pointer)
}

fn openxrextensionwrapper_gd_set_session_create_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetSessionCreateAndGetNextPointer(unsafe{&T(voidptr(inst))})
	next_pointer := unsafe{&voidptr(args[0])}
	*(&i64(ret)) := v_inst.set_session_create_and_get_next_pointer_(next_pointer)
}

fn openxrextensionwrapper_gd_set_swapchain_create_info_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetSwapchainCreateInfoAndGetNextPointer(unsafe{&T(voidptr(inst))})
	next_pointer := unsafe{&voidptr(args[0])}
	*(&i64(ret)) := v_inst.set_swapchain_create_info_and_get_next_pointer_(next_pointer)
}

fn openxrextensionwrapper_gd_set_hand_joint_locations_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetHandJointLocationsAndGetNextPointer(unsafe{&T(voidptr(inst))})
	hand_index := unsafe{&i64(args[0])}
	next_pointer := unsafe{&voidptr(args[1])}
	*(&i64(ret)) := v_inst.set_hand_joint_locations_and_get_next_pointer_(hand_index, next_pointer)
}

fn openxrextensionwrapper_gd_set_projection_views_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetProjectionViewsAndGetNextPointer(unsafe{&T(voidptr(inst))})
	view_index := unsafe{&i64(args[0])}
	next_pointer := unsafe{&voidptr(args[1])}
	*(&i64(ret)) := v_inst.set_projection_views_and_get_next_pointer_(view_index, next_pointer)
}

fn openxrextensionwrapper_gd_set_frame_wait_info_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetFrameWaitInfoAndGetNextPointer(unsafe{&T(voidptr(inst))})
	next_pointer := unsafe{&voidptr(args[0])}
	*(&i64(ret)) := v_inst.set_frame_wait_info_and_get_next_pointer_(next_pointer)
}

fn openxrextensionwrapper_gd_set_frame_end_info_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetFrameEndInfoAndGetNextPointer(unsafe{&T(voidptr(inst))})
	next_pointer := unsafe{&voidptr(args[0])}
	*(&i64(ret)) := v_inst.set_frame_end_info_and_get_next_pointer_(next_pointer)
}

fn openxrextensionwrapper_gd_set_view_locate_info_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetViewLocateInfoAndGetNextPointer(unsafe{&T(voidptr(inst))})
	next_pointer := unsafe{&voidptr(args[0])}
	*(&i64(ret)) := v_inst.set_view_locate_info_and_get_next_pointer_(next_pointer)
}

fn openxrextensionwrapper_gd_set_reference_space_create_info_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetReferenceSpaceCreateInfoAndGetNextPointer(unsafe{&T(voidptr(inst))})
	reference_space_type := unsafe{&i64(args[0])}
	next_pointer := unsafe{&voidptr(args[1])}
	*(&i64(ret)) := v_inst.set_reference_space_create_info_and_get_next_pointer_(reference_space_type, next_pointer)
}

fn openxrextensionwrapper_gd_get_composition_layer_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperGetCompositionLayerCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_composition_layer_count_()
}

fn openxrextensionwrapper_gd_get_composition_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperGetCompositionLayer(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_composition_layer_(index)
}

fn openxrextensionwrapper_gd_get_composition_layer_order[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperGetCompositionLayerOrder(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_composition_layer_order_(index)
}

fn openxrextensionwrapper_gd_get_suggested_tracker_names[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperGetSuggestedTrackerNames(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_suggested_tracker_names_()
}

fn openxrextensionwrapper_gd_on_register_metadata[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnRegisterMetadata(unsafe{&T(voidptr(inst))})
	v_inst.on_register_metadata_()
}

fn openxrextensionwrapper_gd_on_before_instance_created[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnBeforeInstanceCreated(unsafe{&T(voidptr(inst))})
	v_inst.on_before_instance_created_()
}

fn openxrextensionwrapper_gd_on_instance_created[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnInstanceCreated(unsafe{&T(voidptr(inst))})
	instance := unsafe{&i64(args[0])}
	v_inst.on_instance_created_(instance)
}

fn openxrextensionwrapper_gd_on_instance_destroyed[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnInstanceDestroyed(unsafe{&T(voidptr(inst))})
	v_inst.on_instance_destroyed_()
}

fn openxrextensionwrapper_gd_on_session_created[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnSessionCreated(unsafe{&T(voidptr(inst))})
	session := unsafe{&i64(args[0])}
	v_inst.on_session_created_(session)
}

fn openxrextensionwrapper_gd_on_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnProcess(unsafe{&T(voidptr(inst))})
	v_inst.on_process_()
}

fn openxrextensionwrapper_gd_on_pre_render[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnPreRender(unsafe{&T(voidptr(inst))})
	v_inst.on_pre_render_()
}

fn openxrextensionwrapper_gd_on_main_swapchains_created[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnMainSwapchainsCreated(unsafe{&T(voidptr(inst))})
	v_inst.on_main_swapchains_created_()
}

fn openxrextensionwrapper_gd_on_pre_draw_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnPreDrawViewport(unsafe{&T(voidptr(inst))})
	viewport := unsafe{&RID(args[0])}
	v_inst.on_pre_draw_viewport_(viewport)
}

fn openxrextensionwrapper_gd_on_post_draw_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnPostDrawViewport(unsafe{&T(voidptr(inst))})
	viewport := unsafe{&RID(args[0])}
	v_inst.on_post_draw_viewport_(viewport)
}

fn openxrextensionwrapper_gd_on_session_destroyed[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnSessionDestroyed(unsafe{&T(voidptr(inst))})
	v_inst.on_session_destroyed_()
}

fn openxrextensionwrapper_gd_on_state_idle[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateIdle(unsafe{&T(voidptr(inst))})
	v_inst.on_state_idle_()
}

fn openxrextensionwrapper_gd_on_state_ready[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateReady(unsafe{&T(voidptr(inst))})
	v_inst.on_state_ready_()
}

fn openxrextensionwrapper_gd_on_state_synchronized[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateSynchronized(unsafe{&T(voidptr(inst))})
	v_inst.on_state_synchronized_()
}

fn openxrextensionwrapper_gd_on_state_visible[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateVisible(unsafe{&T(voidptr(inst))})
	v_inst.on_state_visible_()
}

fn openxrextensionwrapper_gd_on_state_focused[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateFocused(unsafe{&T(voidptr(inst))})
	v_inst.on_state_focused_()
}

fn openxrextensionwrapper_gd_on_state_stopping[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateStopping(unsafe{&T(voidptr(inst))})
	v_inst.on_state_stopping_()
}

fn openxrextensionwrapper_gd_on_state_loss_pending[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateLossPending(unsafe{&T(voidptr(inst))})
	v_inst.on_state_loss_pending_()
}

fn openxrextensionwrapper_gd_on_state_exiting[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnStateExiting(unsafe{&T(voidptr(inst))})
	v_inst.on_state_exiting_()
}

fn openxrextensionwrapper_gd_on_event_polled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnEventPolled(unsafe{&T(voidptr(inst))})
	event := unsafe{&voidptr(args[0])}
	*(&bool(ret)) := v_inst.on_event_polled_(event)
}

fn openxrextensionwrapper_gd_set_viewport_composition_layer_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetViewportCompositionLayerAndGetNextPointer(unsafe{&T(voidptr(inst))})
	layer := unsafe{&voidptr(args[0])}
	property_values := unsafe{&Dictionary(args[1])}
	next_pointer := unsafe{&voidptr(args[2])}
	*(&i64(ret)) := v_inst.set_viewport_composition_layer_and_get_next_pointer_(layer, property_values, next_pointer)
}

fn openxrextensionwrapper_gd_get_viewport_composition_layer_extension_properties[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperGetViewportCompositionLayerExtensionProperties(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_viewport_composition_layer_extension_properties_()
}

fn openxrextensionwrapper_gd_get_viewport_composition_layer_extension_property_defaults[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperGetViewportCompositionLayerExtensionPropertyDefaults(unsafe{&T(voidptr(inst))})
	*(&Dictionary(ret)) := v_inst.get_viewport_composition_layer_extension_property_defaults_()
}

fn openxrextensionwrapper_gd_on_viewport_composition_layer_destroyed[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperOnViewportCompositionLayerDestroyed(unsafe{&T(voidptr(inst))})
	layer := unsafe{&voidptr(args[0])}
	v_inst.on_viewport_composition_layer_destroyed_(layer)
}

fn openxrextensionwrapper_gd_set_android_surface_swapchain_create_info_and_get_next_pointer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IOpenXRExtensionWrapperSetAndroidSurfaceSwapchainCreateInfoAndGetNextPointer(unsafe{&T(voidptr(inst))})
	property_values := unsafe{&Dictionary(args[0])}
	next_pointer := unsafe{&voidptr(args[1])}
	*(&i64(ret)) := v_inst.set_android_surface_swapchain_create_info_and_get_next_pointer_(property_values, next_pointer)
}

fn packetpeerextension_gd_get_packet[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPacketPeerExtensionGetPacket(unsafe{&T(voidptr(inst))})
	r_buffer := unsafe{&&&u8 (args[0])}
	r_buffer_size := unsafe{&&i32(args[1])}
	*(&GDError(ret)) := v_inst.get_packet_(r_buffer, r_buffer_size)
}

fn packetpeerextension_gd_put_packet[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPacketPeerExtensionPutPacket(unsafe{&T(voidptr(inst))})
	p_buffer := unsafe{&&u8(args[0])}
	p_buffer_size := unsafe{&i64(args[1])}
	*(&GDError(ret)) := v_inst.put_packet_(p_buffer, p_buffer_size)
}

fn packetpeerextension_gd_get_available_packet_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPacketPeerExtensionGetAvailablePacketCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_available_packet_count_()
}

fn packetpeerextension_gd_get_max_packet_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPacketPeerExtensionGetMaxPacketSize(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_max_packet_size_()
}

fn physicalbone3d_gd_integrate_forces[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicalBone3DIntegrateForces(unsafe{&T(voidptr(inst))})
	state := unsafe{&PhysicsDirectBodyState3D(args[0])}
	v_inst.integrate_forces_(state)
}

fn physicsdirectbodystate2dextension_gd_get_total_gravity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetTotalGravity(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_total_gravity_()
}

fn physicsdirectbodystate2dextension_gd_get_total_linear_damp[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetTotalLinearDamp(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_total_linear_damp_()
}

fn physicsdirectbodystate2dextension_gd_get_total_angular_damp[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetTotalAngularDamp(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_total_angular_damp_()
}

fn physicsdirectbodystate2dextension_gd_get_center_of_mass[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetCenterOfMass(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_center_of_mass_()
}

fn physicsdirectbodystate2dextension_gd_get_center_of_mass_local[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetCenterOfMassLocal(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_center_of_mass_local_()
}

fn physicsdirectbodystate2dextension_gd_get_inverse_mass[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetInverseMass(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_inverse_mass_()
}

fn physicsdirectbodystate2dextension_gd_get_inverse_inertia[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetInverseInertia(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_inverse_inertia_()
}

fn physicsdirectbodystate2dextension_gd_set_linear_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionSetLinearVelocity(unsafe{&T(voidptr(inst))})
	velocity := unsafe{&Vector2(args[0])}
	v_inst.set_linear_velocity_(velocity)
}

fn physicsdirectbodystate2dextension_gd_get_linear_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetLinearVelocity(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_linear_velocity_()
}

fn physicsdirectbodystate2dextension_gd_set_angular_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionSetAngularVelocity(unsafe{&T(voidptr(inst))})
	velocity := unsafe{&f64(args[0])}
	v_inst.set_angular_velocity_(velocity)
}

fn physicsdirectbodystate2dextension_gd_get_angular_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetAngularVelocity(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_angular_velocity_()
}

fn physicsdirectbodystate2dextension_gd_set_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionSetTransform(unsafe{&T(voidptr(inst))})
	transform := unsafe{&Transform2D(args[0])}
	v_inst.set_transform_(transform)
}

fn physicsdirectbodystate2dextension_gd_get_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetTransform(unsafe{&T(voidptr(inst))})
	*(&Transform2D(ret)) := v_inst.get_transform_()
}

fn physicsdirectbodystate2dextension_gd_get_velocity_at_local_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetVelocityAtLocalPosition(unsafe{&T(voidptr(inst))})
	local_position := unsafe{&Vector2(args[0])}
	*(&Vector2(ret)) := v_inst.get_velocity_at_local_position_(local_position)
}

fn physicsdirectbodystate2dextension_gd_apply_central_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionApplyCentralImpulse(unsafe{&T(voidptr(inst))})
	impulse := unsafe{&Vector2(args[0])}
	v_inst.apply_central_impulse_(impulse)
}

fn physicsdirectbodystate2dextension_gd_apply_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionApplyImpulse(unsafe{&T(voidptr(inst))})
	impulse := unsafe{&Vector2(args[0])}
	position := unsafe{&Vector2(args[1])}
	v_inst.apply_impulse_(impulse, position)
}

fn physicsdirectbodystate2dextension_gd_apply_torque_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionApplyTorqueImpulse(unsafe{&T(voidptr(inst))})
	impulse := unsafe{&f64(args[0])}
	v_inst.apply_torque_impulse_(impulse)
}

fn physicsdirectbodystate2dextension_gd_apply_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionApplyCentralForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector2(args[0])}
	v_inst.apply_central_force_(force)
}

fn physicsdirectbodystate2dextension_gd_apply_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionApplyForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector2(args[0])}
	position := unsafe{&Vector2(args[1])}
	v_inst.apply_force_(force, position)
}

fn physicsdirectbodystate2dextension_gd_apply_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionApplyTorque(unsafe{&T(voidptr(inst))})
	torque := unsafe{&f64(args[0])}
	v_inst.apply_torque_(torque)
}

fn physicsdirectbodystate2dextension_gd_add_constant_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionAddConstantCentralForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector2(args[0])}
	v_inst.add_constant_central_force_(force)
}

fn physicsdirectbodystate2dextension_gd_add_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionAddConstantForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector2(args[0])}
	position := unsafe{&Vector2(args[1])}
	v_inst.add_constant_force_(force, position)
}

fn physicsdirectbodystate2dextension_gd_add_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionAddConstantTorque(unsafe{&T(voidptr(inst))})
	torque := unsafe{&f64(args[0])}
	v_inst.add_constant_torque_(torque)
}

fn physicsdirectbodystate2dextension_gd_set_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionSetConstantForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector2(args[0])}
	v_inst.set_constant_force_(force)
}

fn physicsdirectbodystate2dextension_gd_get_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetConstantForce(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_constant_force_()
}

fn physicsdirectbodystate2dextension_gd_set_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionSetConstantTorque(unsafe{&T(voidptr(inst))})
	torque := unsafe{&f64(args[0])}
	v_inst.set_constant_torque_(torque)
}

fn physicsdirectbodystate2dextension_gd_get_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetConstantTorque(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_constant_torque_()
}

fn physicsdirectbodystate2dextension_gd_set_sleep_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionSetSleepState(unsafe{&T(voidptr(inst))})
	enabled := unsafe{&bool(args[0])}
	v_inst.set_sleep_state_(enabled)
}

fn physicsdirectbodystate2dextension_gd_is_sleeping[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionIsSleeping(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_sleeping_()
}

fn physicsdirectbodystate2dextension_gd_get_contact_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_contact_count_()
}

fn physicsdirectbodystate2dextension_gd_get_contact_local_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactLocalPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector2(ret)) := v_inst.get_contact_local_position_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_local_normal[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactLocalNormal(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector2(ret)) := v_inst.get_contact_local_normal_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_local_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactLocalShape(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_contact_local_shape_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_local_velocity_at_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactLocalVelocityAtPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector2(ret)) := v_inst.get_contact_local_velocity_at_position_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_collider[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactCollider(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&RID(ret)) := v_inst.get_contact_collider_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_collider_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactColliderPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector2(ret)) := v_inst.get_contact_collider_position_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_collider_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactColliderId(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_contact_collider_id_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_collider_object[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactColliderObject(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Object(ret)) := v_inst.get_contact_collider_object_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_collider_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactColliderShape(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_contact_collider_shape_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_collider_velocity_at_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactColliderVelocityAtPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector2(ret)) := v_inst.get_contact_collider_velocity_at_position_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_contact_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetContactImpulse(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector2(ret)) := v_inst.get_contact_impulse_(contact_idx)
}

fn physicsdirectbodystate2dextension_gd_get_step[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetStep(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_step_()
}

fn physicsdirectbodystate2dextension_gd_integrate_forces[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionIntegrateForces(unsafe{&T(voidptr(inst))})
	v_inst.integrate_forces_()
}

fn physicsdirectbodystate2dextension_gd_get_space_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState2DExtensionGetSpaceState(unsafe{&T(voidptr(inst))})
	*(&PhysicsDirectSpaceState2D(ret)) := v_inst.get_space_state_()
}

fn physicsdirectbodystate3dextension_gd_get_total_gravity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetTotalGravity(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_total_gravity_()
}

fn physicsdirectbodystate3dextension_gd_get_total_linear_damp[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetTotalLinearDamp(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_total_linear_damp_()
}

fn physicsdirectbodystate3dextension_gd_get_total_angular_damp[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetTotalAngularDamp(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_total_angular_damp_()
}

fn physicsdirectbodystate3dextension_gd_get_center_of_mass[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetCenterOfMass(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_center_of_mass_()
}

fn physicsdirectbodystate3dextension_gd_get_center_of_mass_local[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetCenterOfMassLocal(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_center_of_mass_local_()
}

fn physicsdirectbodystate3dextension_gd_get_principal_inertia_axes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetPrincipalInertiaAxes(unsafe{&T(voidptr(inst))})
	*(&Basis(ret)) := v_inst.get_principal_inertia_axes_()
}

fn physicsdirectbodystate3dextension_gd_get_inverse_mass[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetInverseMass(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_inverse_mass_()
}

fn physicsdirectbodystate3dextension_gd_get_inverse_inertia[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetInverseInertia(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_inverse_inertia_()
}

fn physicsdirectbodystate3dextension_gd_get_inverse_inertia_tensor[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetInverseInertiaTensor(unsafe{&T(voidptr(inst))})
	*(&Basis(ret)) := v_inst.get_inverse_inertia_tensor_()
}

fn physicsdirectbodystate3dextension_gd_set_linear_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionSetLinearVelocity(unsafe{&T(voidptr(inst))})
	velocity := unsafe{&Vector3(args[0])}
	v_inst.set_linear_velocity_(velocity)
}

fn physicsdirectbodystate3dextension_gd_get_linear_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetLinearVelocity(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_linear_velocity_()
}

fn physicsdirectbodystate3dextension_gd_set_angular_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionSetAngularVelocity(unsafe{&T(voidptr(inst))})
	velocity := unsafe{&Vector3(args[0])}
	v_inst.set_angular_velocity_(velocity)
}

fn physicsdirectbodystate3dextension_gd_get_angular_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetAngularVelocity(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_angular_velocity_()
}

fn physicsdirectbodystate3dextension_gd_set_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionSetTransform(unsafe{&T(voidptr(inst))})
	transform := unsafe{&Transform3D(args[0])}
	v_inst.set_transform_(transform)
}

fn physicsdirectbodystate3dextension_gd_get_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetTransform(unsafe{&T(voidptr(inst))})
	*(&Transform3D(ret)) := v_inst.get_transform_()
}

fn physicsdirectbodystate3dextension_gd_get_velocity_at_local_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetVelocityAtLocalPosition(unsafe{&T(voidptr(inst))})
	local_position := unsafe{&Vector3(args[0])}
	*(&Vector3(ret)) := v_inst.get_velocity_at_local_position_(local_position)
}

fn physicsdirectbodystate3dextension_gd_apply_central_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionApplyCentralImpulse(unsafe{&T(voidptr(inst))})
	impulse := unsafe{&Vector3(args[0])}
	v_inst.apply_central_impulse_(impulse)
}

fn physicsdirectbodystate3dextension_gd_apply_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionApplyImpulse(unsafe{&T(voidptr(inst))})
	impulse := unsafe{&Vector3(args[0])}
	position := unsafe{&Vector3(args[1])}
	v_inst.apply_impulse_(impulse, position)
}

fn physicsdirectbodystate3dextension_gd_apply_torque_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionApplyTorqueImpulse(unsafe{&T(voidptr(inst))})
	impulse := unsafe{&Vector3(args[0])}
	v_inst.apply_torque_impulse_(impulse)
}

fn physicsdirectbodystate3dextension_gd_apply_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionApplyCentralForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector3(args[0])}
	v_inst.apply_central_force_(force)
}

fn physicsdirectbodystate3dextension_gd_apply_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionApplyForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector3(args[0])}
	position := unsafe{&Vector3(args[1])}
	v_inst.apply_force_(force, position)
}

fn physicsdirectbodystate3dextension_gd_apply_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionApplyTorque(unsafe{&T(voidptr(inst))})
	torque := unsafe{&Vector3(args[0])}
	v_inst.apply_torque_(torque)
}

fn physicsdirectbodystate3dextension_gd_add_constant_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionAddConstantCentralForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector3(args[0])}
	v_inst.add_constant_central_force_(force)
}

fn physicsdirectbodystate3dextension_gd_add_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionAddConstantForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector3(args[0])}
	position := unsafe{&Vector3(args[1])}
	v_inst.add_constant_force_(force, position)
}

fn physicsdirectbodystate3dextension_gd_add_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionAddConstantTorque(unsafe{&T(voidptr(inst))})
	torque := unsafe{&Vector3(args[0])}
	v_inst.add_constant_torque_(torque)
}

fn physicsdirectbodystate3dextension_gd_set_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionSetConstantForce(unsafe{&T(voidptr(inst))})
	force := unsafe{&Vector3(args[0])}
	v_inst.set_constant_force_(force)
}

fn physicsdirectbodystate3dextension_gd_get_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetConstantForce(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_constant_force_()
}

fn physicsdirectbodystate3dextension_gd_set_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionSetConstantTorque(unsafe{&T(voidptr(inst))})
	torque := unsafe{&Vector3(args[0])}
	v_inst.set_constant_torque_(torque)
}

fn physicsdirectbodystate3dextension_gd_get_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetConstantTorque(unsafe{&T(voidptr(inst))})
	*(&Vector3(ret)) := v_inst.get_constant_torque_()
}

fn physicsdirectbodystate3dextension_gd_set_sleep_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionSetSleepState(unsafe{&T(voidptr(inst))})
	enabled := unsafe{&bool(args[0])}
	v_inst.set_sleep_state_(enabled)
}

fn physicsdirectbodystate3dextension_gd_is_sleeping[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionIsSleeping(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_sleeping_()
}

fn physicsdirectbodystate3dextension_gd_get_contact_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_contact_count_()
}

fn physicsdirectbodystate3dextension_gd_get_contact_local_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactLocalPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector3(ret)) := v_inst.get_contact_local_position_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_local_normal[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactLocalNormal(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector3(ret)) := v_inst.get_contact_local_normal_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactImpulse(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector3(ret)) := v_inst.get_contact_impulse_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_local_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactLocalShape(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_contact_local_shape_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_local_velocity_at_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactLocalVelocityAtPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector3(ret)) := v_inst.get_contact_local_velocity_at_position_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_collider[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactCollider(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&RID(ret)) := v_inst.get_contact_collider_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_collider_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactColliderPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector3(ret)) := v_inst.get_contact_collider_position_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_collider_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactColliderId(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_contact_collider_id_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_collider_object[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactColliderObject(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Object(ret)) := v_inst.get_contact_collider_object_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_collider_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactColliderShape(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_contact_collider_shape_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_contact_collider_velocity_at_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetContactColliderVelocityAtPosition(unsafe{&T(voidptr(inst))})
	contact_idx := unsafe{&i64(args[0])}
	*(&Vector3(ret)) := v_inst.get_contact_collider_velocity_at_position_(contact_idx)
}

fn physicsdirectbodystate3dextension_gd_get_step[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetStep(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_step_()
}

fn physicsdirectbodystate3dextension_gd_integrate_forces[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionIntegrateForces(unsafe{&T(voidptr(inst))})
	v_inst.integrate_forces_()
}

fn physicsdirectbodystate3dextension_gd_get_space_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectBodyState3DExtensionGetSpaceState(unsafe{&T(voidptr(inst))})
	*(&PhysicsDirectSpaceState3D(ret)) := v_inst.get_space_state_()
}

fn physicsdirectspacestate2dextension_gd_intersect_ray[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState2DExtensionIntersectRay(unsafe{&T(voidptr(inst))})
	from := unsafe{&Vector2(args[0])}
	to := unsafe{&Vector2(args[1])}
	collision_mask := unsafe{&i64(args[2])}
	collide_with_bodies := unsafe{&bool(args[3])}
	collide_with_areas := unsafe{&bool(args[4])}
	hit_from_inside := unsafe{&bool(args[5])}
	gd_result := unsafe{&&PhysicsServer2DExtensionRayResult(args[6])}
	*(&bool(ret)) := v_inst.intersect_ray_(from, to, collision_mask, collide_with_bodies, collide_with_areas, hit_from_inside, gd_result)
}

fn physicsdirectspacestate2dextension_gd_intersect_point[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState2DExtensionIntersectPoint(unsafe{&T(voidptr(inst))})
	position := unsafe{&Vector2(args[0])}
	canvas_instance_id := unsafe{&i64(args[1])}
	collision_mask := unsafe{&i64(args[2])}
	collide_with_bodies := unsafe{&bool(args[3])}
	collide_with_areas := unsafe{&bool(args[4])}
	results := unsafe{&&PhysicsServer2DExtensionShapeResult(args[5])}
	max_results := unsafe{&i64(args[6])}
	*(&i64(ret)) := v_inst.intersect_point_(position, canvas_instance_id, collision_mask, collide_with_bodies, collide_with_areas, results, max_results)
}

fn physicsdirectspacestate2dextension_gd_intersect_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState2DExtensionIntersectShape(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform2D(args[1])}
	motion := unsafe{&Vector2(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	gd_result := unsafe{&&PhysicsServer2DExtensionShapeResult(args[7])}
	max_results := unsafe{&i64(args[8])}
	*(&i64(ret)) := v_inst.intersect_shape_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, gd_result, max_results)
}

fn physicsdirectspacestate2dextension_gd_cast_motion[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState2DExtensionCastMotion(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform2D(args[1])}
	motion := unsafe{&Vector2(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	closest_safe := unsafe{&&f64(args[7])}
	closest_unsafe := unsafe{&&f64(args[8])}
	*(&bool(ret)) := v_inst.cast_motion_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, closest_safe, closest_unsafe)
}

fn physicsdirectspacestate2dextension_gd_collide_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState2DExtensionCollideShape(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform2D(args[1])}
	motion := unsafe{&Vector2(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	results := unsafe{&voidptr(args[7])}
	max_results := unsafe{&i64(args[8])}
	result_count := unsafe{&&i32(args[9])}
	*(&bool(ret)) := v_inst.collide_shape_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, results, max_results, result_count)
}

fn physicsdirectspacestate2dextension_gd_rest_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState2DExtensionRestInfo(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform2D(args[1])}
	motion := unsafe{&Vector2(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	rest_info := unsafe{&&PhysicsServer2DExtensionShapeRestInfo(args[7])}
	*(&bool(ret)) := v_inst.rest_info_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, rest_info)
}

fn physicsdirectspacestate3dextension_gd_intersect_ray[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState3DExtensionIntersectRay(unsafe{&T(voidptr(inst))})
	from := unsafe{&Vector3(args[0])}
	to := unsafe{&Vector3(args[1])}
	collision_mask := unsafe{&i64(args[2])}
	collide_with_bodies := unsafe{&bool(args[3])}
	collide_with_areas := unsafe{&bool(args[4])}
	hit_from_inside := unsafe{&bool(args[5])}
	hit_back_faces := unsafe{&bool(args[6])}
	pick_ray := unsafe{&bool(args[7])}
	gd_result := unsafe{&&PhysicsServer3DExtensionRayResult(args[8])}
	*(&bool(ret)) := v_inst.intersect_ray_(from, to, collision_mask, collide_with_bodies, collide_with_areas, hit_from_inside, hit_back_faces, pick_ray, gd_result)
}

fn physicsdirectspacestate3dextension_gd_intersect_point[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState3DExtensionIntersectPoint(unsafe{&T(voidptr(inst))})
	position := unsafe{&Vector3(args[0])}
	collision_mask := unsafe{&i64(args[1])}
	collide_with_bodies := unsafe{&bool(args[2])}
	collide_with_areas := unsafe{&bool(args[3])}
	results := unsafe{&&PhysicsServer3DExtensionShapeResult(args[4])}
	max_results := unsafe{&i64(args[5])}
	*(&i64(ret)) := v_inst.intersect_point_(position, collision_mask, collide_with_bodies, collide_with_areas, results, max_results)
}

fn physicsdirectspacestate3dextension_gd_intersect_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState3DExtensionIntersectShape(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform3D(args[1])}
	motion := unsafe{&Vector3(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	result_count := unsafe{&&PhysicsServer3DExtensionShapeResult(args[7])}
	max_results := unsafe{&i64(args[8])}
	*(&i64(ret)) := v_inst.intersect_shape_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, result_count, max_results)
}

fn physicsdirectspacestate3dextension_gd_cast_motion[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState3DExtensionCastMotion(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform3D(args[1])}
	motion := unsafe{&Vector3(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	closest_safe := unsafe{&&f64(args[7])}
	closest_unsafe := unsafe{&&f64(args[8])}
	info := unsafe{&&PhysicsServer3DExtensionShapeRestInfo(args[9])}
	*(&bool(ret)) := v_inst.cast_motion_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, closest_safe, closest_unsafe, info)
}

fn physicsdirectspacestate3dextension_gd_collide_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState3DExtensionCollideShape(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform3D(args[1])}
	motion := unsafe{&Vector3(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	results := unsafe{&voidptr(args[7])}
	max_results := unsafe{&i64(args[8])}
	result_count := unsafe{&&i32(args[9])}
	*(&bool(ret)) := v_inst.collide_shape_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, results, max_results, result_count)
}

fn physicsdirectspacestate3dextension_gd_rest_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState3DExtensionRestInfo(unsafe{&T(voidptr(inst))})
	shape_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform3D(args[1])}
	motion := unsafe{&Vector3(args[2])}
	margin := unsafe{&f64(args[3])}
	collision_mask := unsafe{&i64(args[4])}
	collide_with_bodies := unsafe{&bool(args[5])}
	collide_with_areas := unsafe{&bool(args[6])}
	rest_info := unsafe{&&PhysicsServer3DExtensionShapeRestInfo(args[7])}
	*(&bool(ret)) := v_inst.rest_info_(shape_rid, transform, motion, margin, collision_mask, collide_with_bodies, collide_with_areas, rest_info)
}

fn physicsdirectspacestate3dextension_gd_get_closest_point_to_object_volume[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsDirectSpaceState3DExtensionGetClosestPointToObjectVolume(unsafe{&T(voidptr(inst))})
	object := unsafe{&RID(args[0])}
	point := unsafe{&Vector3(args[1])}
	*(&Vector3(ret)) := v_inst.get_closest_point_to_object_volume_(object, point)
}

fn physicsserver2dextension_gd_world_boundary_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionWorldBoundaryShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.world_boundary_shape_create_()
}

fn physicsserver2dextension_gd_separation_ray_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSeparationRayShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.separation_ray_shape_create_()
}

fn physicsserver2dextension_gd_segment_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSegmentShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.segment_shape_create_()
}

fn physicsserver2dextension_gd_circle_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionCircleShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.circle_shape_create_()
}

fn physicsserver2dextension_gd_rectangle_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionRectangleShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.rectangle_shape_create_()
}

fn physicsserver2dextension_gd_capsule_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionCapsuleShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.capsule_shape_create_()
}

fn physicsserver2dextension_gd_convex_polygon_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionConvexPolygonShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.convex_polygon_shape_create_()
}

fn physicsserver2dextension_gd_concave_polygon_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionConcavePolygonShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.concave_polygon_shape_create_()
}

fn physicsserver2dextension_gd_shape_set_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionShapeSetData(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	data := unsafe{&Variant(args[1])}
	v_inst.shape_set_data_(shape, data)
}

fn physicsserver2dextension_gd_shape_set_custom_solver_bias[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionShapeSetCustomSolverBias(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	bias := unsafe{&f64(args[1])}
	v_inst.shape_set_custom_solver_bias_(shape, bias)
}

fn physicsserver2dextension_gd_shape_get_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionShapeGetType(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	*(&PhysicsServer2DShapeType(ret)) := v_inst.shape_get_type_(shape)
}

fn physicsserver2dextension_gd_shape_get_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionShapeGetData(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	*(&Variant(ret)) := v_inst.shape_get_data_(shape)
}

fn physicsserver2dextension_gd_shape_get_custom_solver_bias[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionShapeGetCustomSolverBias(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shape_get_custom_solver_bias_(shape)
}

fn physicsserver2dextension_gd_shape_collide[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionShapeCollide(unsafe{&T(voidptr(inst))})
	shape_a := unsafe{&RID(args[0])}
	xform_a := unsafe{&Transform2D(args[1])}
	motion_a := unsafe{&Vector2(args[2])}
	shape_b := unsafe{&RID(args[3])}
	xform_b := unsafe{&Transform2D(args[4])}
	motion_b := unsafe{&Vector2(args[5])}
	results := unsafe{&voidptr(args[6])}
	result_max := unsafe{&i64(args[7])}
	result_count := unsafe{&&i32(args[8])}
	*(&bool(ret)) := v_inst.shape_collide_(shape_a, xform_a, motion_a, shape_b, xform_b, motion_b, results, result_max, result_count)
}

fn physicsserver2dextension_gd_space_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.space_create_()
}

fn physicsserver2dextension_gd_space_set_active[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceSetActive(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	active := unsafe{&bool(args[1])}
	v_inst.space_set_active_(space, active)
}

fn physicsserver2dextension_gd_space_is_active[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceIsActive(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.space_is_active_(space)
}

fn physicsserver2dextension_gd_space_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceSetParam(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DSpaceParameter(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.space_set_param_(space, param, value)
}

fn physicsserver2dextension_gd_space_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceGetParam(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DSpaceParameter(args[1])}
	*(&f64(ret)) := v_inst.space_get_param_(space, param)
}

fn physicsserver2dextension_gd_space_get_direct_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceGetDirectState(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&PhysicsDirectSpaceState2D(ret)) := v_inst.space_get_direct_state_(space)
}

fn physicsserver2dextension_gd_space_set_debug_contacts[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceSetDebugContacts(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	max_contacts := unsafe{&i64(args[1])}
	v_inst.space_set_debug_contacts_(space, max_contacts)
}

fn physicsserver2dextension_gd_space_get_contacts[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceGetContacts(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&PackedVector2Array(ret)) := v_inst.space_get_contacts_(space)
}

fn physicsserver2dextension_gd_space_get_contact_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSpaceGetContactCount(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.space_get_contact_count_(space)
}

fn physicsserver2dextension_gd_area_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.area_create_()
}

fn physicsserver2dextension_gd_area_set_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetSpace(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	space := unsafe{&RID(args[1])}
	v_inst.area_set_space_(area, space)
}

fn physicsserver2dextension_gd_area_get_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetSpace(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&RID(ret)) := v_inst.area_get_space_(area)
}

fn physicsserver2dextension_gd_area_add_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaAddShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape := unsafe{&RID(args[1])}
	transform := unsafe{&Transform2D(args[2])}
	disabled := unsafe{&bool(args[3])}
	v_inst.area_add_shape_(area, shape, transform, disabled)
}

fn physicsserver2dextension_gd_area_set_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	shape := unsafe{&RID(args[2])}
	v_inst.area_set_shape_(area, shape_idx, shape)
}

fn physicsserver2dextension_gd_area_set_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetShapeTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	transform := unsafe{&Transform2D(args[2])}
	v_inst.area_set_shape_transform_(area, shape_idx, transform)
}

fn physicsserver2dextension_gd_area_set_shape_disabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetShapeDisabled(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	disabled := unsafe{&bool(args[2])}
	v_inst.area_set_shape_disabled_(area, shape_idx, disabled)
}

fn physicsserver2dextension_gd_area_get_shape_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetShapeCount(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_shape_count_(area)
}

fn physicsserver2dextension_gd_area_get_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&RID(ret)) := v_inst.area_get_shape_(area, shape_idx)
}

fn physicsserver2dextension_gd_area_get_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetShapeTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&Transform2D(ret)) := v_inst.area_get_shape_transform_(area, shape_idx)
}

fn physicsserver2dextension_gd_area_remove_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaRemoveShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	v_inst.area_remove_shape_(area, shape_idx)
}

fn physicsserver2dextension_gd_area_clear_shapes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaClearShapes(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	v_inst.area_clear_shapes_(area)
}

fn physicsserver2dextension_gd_area_attach_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaAttachObjectInstanceId(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	id := unsafe{&i64(args[1])}
	v_inst.area_attach_object_instance_id_(area, id)
}

fn physicsserver2dextension_gd_area_get_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetObjectInstanceId(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_object_instance_id_(area)
}

fn physicsserver2dextension_gd_area_attach_canvas_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaAttachCanvasInstanceId(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	id := unsafe{&i64(args[1])}
	v_inst.area_attach_canvas_instance_id_(area, id)
}

fn physicsserver2dextension_gd_area_get_canvas_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetCanvasInstanceId(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_canvas_instance_id_(area)
}

fn physicsserver2dextension_gd_area_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetParam(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DAreaParameter(args[1])}
	value := unsafe{&Variant(args[2])}
	v_inst.area_set_param_(area, param, value)
}

fn physicsserver2dextension_gd_area_set_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	transform := unsafe{&Transform2D(args[1])}
	v_inst.area_set_transform_(area, transform)
}

fn physicsserver2dextension_gd_area_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetParam(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DAreaParameter(args[1])}
	*(&Variant(ret)) := v_inst.area_get_param_(area, param)
}

fn physicsserver2dextension_gd_area_get_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&Transform2D(ret)) := v_inst.area_get_transform_(area)
}

fn physicsserver2dextension_gd_area_set_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetCollisionLayer(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	layer := unsafe{&i64(args[1])}
	v_inst.area_set_collision_layer_(area, layer)
}

fn physicsserver2dextension_gd_area_get_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetCollisionLayer(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_collision_layer_(area)
}

fn physicsserver2dextension_gd_area_set_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetCollisionMask(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	mask := unsafe{&i64(args[1])}
	v_inst.area_set_collision_mask_(area, mask)
}

fn physicsserver2dextension_gd_area_get_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaGetCollisionMask(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_collision_mask_(area)
}

fn physicsserver2dextension_gd_area_set_monitorable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetMonitorable(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	monitorable := unsafe{&bool(args[1])}
	v_inst.area_set_monitorable_(area, monitorable)
}

fn physicsserver2dextension_gd_area_set_pickable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetPickable(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	pickable := unsafe{&bool(args[1])}
	v_inst.area_set_pickable_(area, pickable)
}

fn physicsserver2dextension_gd_area_set_monitor_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetMonitorCallback(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	callback := unsafe{&Callable(args[1])}
	v_inst.area_set_monitor_callback_(area, callback)
}

fn physicsserver2dextension_gd_area_set_area_monitor_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionAreaSetAreaMonitorCallback(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	callback := unsafe{&Callable(args[1])}
	v_inst.area_set_area_monitor_callback_(area, callback)
}

fn physicsserver2dextension_gd_body_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.body_create_()
}

fn physicsserver2dextension_gd_body_set_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetSpace(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	space := unsafe{&RID(args[1])}
	v_inst.body_set_space_(body, space)
}

fn physicsserver2dextension_gd_body_get_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetSpace(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&RID(ret)) := v_inst.body_get_space_(body)
}

fn physicsserver2dextension_gd_body_set_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetMode(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	mode := unsafe{&PhysicsServer2DBodyMode(args[1])}
	v_inst.body_set_mode_(body, mode)
}

fn physicsserver2dextension_gd_body_get_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetMode(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&PhysicsServer2DBodyMode(ret)) := v_inst.body_get_mode_(body)
}

fn physicsserver2dextension_gd_body_add_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyAddShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape := unsafe{&RID(args[1])}
	transform := unsafe{&Transform2D(args[2])}
	disabled := unsafe{&bool(args[3])}
	v_inst.body_add_shape_(body, shape, transform, disabled)
}

fn physicsserver2dextension_gd_body_set_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	shape := unsafe{&RID(args[2])}
	v_inst.body_set_shape_(body, shape_idx, shape)
}

fn physicsserver2dextension_gd_body_set_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetShapeTransform(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	transform := unsafe{&Transform2D(args[2])}
	v_inst.body_set_shape_transform_(body, shape_idx, transform)
}

fn physicsserver2dextension_gd_body_get_shape_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetShapeCount(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_shape_count_(body)
}

fn physicsserver2dextension_gd_body_get_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&RID(ret)) := v_inst.body_get_shape_(body, shape_idx)
}

fn physicsserver2dextension_gd_body_get_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetShapeTransform(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&Transform2D(ret)) := v_inst.body_get_shape_transform_(body, shape_idx)
}

fn physicsserver2dextension_gd_body_set_shape_disabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetShapeDisabled(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	disabled := unsafe{&bool(args[2])}
	v_inst.body_set_shape_disabled_(body, shape_idx, disabled)
}

fn physicsserver2dextension_gd_body_set_shape_as_one_way_collision[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetShapeAsOneWayCollision(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	enable := unsafe{&bool(args[2])}
	margin := unsafe{&f64(args[3])}
	v_inst.body_set_shape_as_one_way_collision_(body, shape_idx, enable, margin)
}

fn physicsserver2dextension_gd_body_remove_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyRemoveShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	v_inst.body_remove_shape_(body, shape_idx)
}

fn physicsserver2dextension_gd_body_clear_shapes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyClearShapes(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	v_inst.body_clear_shapes_(body)
}

fn physicsserver2dextension_gd_body_attach_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyAttachObjectInstanceId(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	id := unsafe{&i64(args[1])}
	v_inst.body_attach_object_instance_id_(body, id)
}

fn physicsserver2dextension_gd_body_get_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetObjectInstanceId(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_object_instance_id_(body)
}

fn physicsserver2dextension_gd_body_attach_canvas_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyAttachCanvasInstanceId(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	id := unsafe{&i64(args[1])}
	v_inst.body_attach_canvas_instance_id_(body, id)
}

fn physicsserver2dextension_gd_body_get_canvas_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetCanvasInstanceId(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_canvas_instance_id_(body)
}

fn physicsserver2dextension_gd_body_set_continuous_collision_detection_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetContinuousCollisionDetectionMode(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	mode := unsafe{&PhysicsServer2DCCDMode(args[1])}
	v_inst.body_set_continuous_collision_detection_mode_(body, mode)
}

fn physicsserver2dextension_gd_body_get_continuous_collision_detection_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetContinuousCollisionDetectionMode(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&PhysicsServer2DCCDMode(ret)) := v_inst.body_get_continuous_collision_detection_mode_(body)
}

fn physicsserver2dextension_gd_body_set_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetCollisionLayer(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	layer := unsafe{&i64(args[1])}
	v_inst.body_set_collision_layer_(body, layer)
}

fn physicsserver2dextension_gd_body_get_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetCollisionLayer(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_collision_layer_(body)
}

fn physicsserver2dextension_gd_body_set_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetCollisionMask(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	mask := unsafe{&i64(args[1])}
	v_inst.body_set_collision_mask_(body, mask)
}

fn physicsserver2dextension_gd_body_get_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetCollisionMask(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_collision_mask_(body)
}

fn physicsserver2dextension_gd_body_set_collision_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetCollisionPriority(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	priority := unsafe{&f64(args[1])}
	v_inst.body_set_collision_priority_(body, priority)
}

fn physicsserver2dextension_gd_body_get_collision_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetCollisionPriority(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.body_get_collision_priority_(body)
}

fn physicsserver2dextension_gd_body_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetParam(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DBodyParameter(args[1])}
	value := unsafe{&Variant(args[2])}
	v_inst.body_set_param_(body, param, value)
}

fn physicsserver2dextension_gd_body_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetParam(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DBodyParameter(args[1])}
	*(&Variant(ret)) := v_inst.body_get_param_(body, param)
}

fn physicsserver2dextension_gd_body_reset_mass_properties[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyResetMassProperties(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	v_inst.body_reset_mass_properties_(body)
}

fn physicsserver2dextension_gd_body_set_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	state := unsafe{&PhysicsServer2DBodyState(args[1])}
	value := unsafe{&Variant(args[2])}
	v_inst.body_set_state_(body, state, value)
}

fn physicsserver2dextension_gd_body_get_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	state := unsafe{&PhysicsServer2DBodyState(args[1])}
	*(&Variant(ret)) := v_inst.body_get_state_(body, state)
}

fn physicsserver2dextension_gd_body_apply_central_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyApplyCentralImpulse(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	impulse := unsafe{&Vector2(args[1])}
	v_inst.body_apply_central_impulse_(body, impulse)
}

fn physicsserver2dextension_gd_body_apply_torque_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyApplyTorqueImpulse(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	impulse := unsafe{&f64(args[1])}
	v_inst.body_apply_torque_impulse_(body, impulse)
}

fn physicsserver2dextension_gd_body_apply_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyApplyImpulse(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	impulse := unsafe{&Vector2(args[1])}
	position := unsafe{&Vector2(args[2])}
	v_inst.body_apply_impulse_(body, impulse, position)
}

fn physicsserver2dextension_gd_body_apply_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyApplyCentralForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector2(args[1])}
	v_inst.body_apply_central_force_(body, force)
}

fn physicsserver2dextension_gd_body_apply_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyApplyForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector2(args[1])}
	position := unsafe{&Vector2(args[2])}
	v_inst.body_apply_force_(body, force, position)
}

fn physicsserver2dextension_gd_body_apply_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyApplyTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	torque := unsafe{&f64(args[1])}
	v_inst.body_apply_torque_(body, torque)
}

fn physicsserver2dextension_gd_body_add_constant_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyAddConstantCentralForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector2(args[1])}
	v_inst.body_add_constant_central_force_(body, force)
}

fn physicsserver2dextension_gd_body_add_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyAddConstantForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector2(args[1])}
	position := unsafe{&Vector2(args[2])}
	v_inst.body_add_constant_force_(body, force, position)
}

fn physicsserver2dextension_gd_body_add_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyAddConstantTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	torque := unsafe{&f64(args[1])}
	v_inst.body_add_constant_torque_(body, torque)
}

fn physicsserver2dextension_gd_body_set_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetConstantForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector2(args[1])}
	v_inst.body_set_constant_force_(body, force)
}

fn physicsserver2dextension_gd_body_get_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetConstantForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&Vector2(ret)) := v_inst.body_get_constant_force_(body)
}

fn physicsserver2dextension_gd_body_set_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetConstantTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	torque := unsafe{&f64(args[1])}
	v_inst.body_set_constant_torque_(body, torque)
}

fn physicsserver2dextension_gd_body_get_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetConstantTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.body_get_constant_torque_(body)
}

fn physicsserver2dextension_gd_body_set_axis_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetAxisVelocity(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	axis_velocity := unsafe{&Vector2(args[1])}
	v_inst.body_set_axis_velocity_(body, axis_velocity)
}

fn physicsserver2dextension_gd_body_add_collision_exception[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyAddCollisionException(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	excepted_body := unsafe{&RID(args[1])}
	v_inst.body_add_collision_exception_(body, excepted_body)
}

fn physicsserver2dextension_gd_body_remove_collision_exception[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyRemoveCollisionException(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	excepted_body := unsafe{&RID(args[1])}
	v_inst.body_remove_collision_exception_(body, excepted_body)
}

fn physicsserver2dextension_gd_body_get_collision_exceptions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetCollisionExceptions(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&Array(ret)) := v_inst.body_get_collision_exceptions_(body)
}

fn physicsserver2dextension_gd_body_set_max_contacts_reported[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetMaxContactsReported(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	amount := unsafe{&i64(args[1])}
	v_inst.body_set_max_contacts_reported_(body, amount)
}

fn physicsserver2dextension_gd_body_get_max_contacts_reported[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetMaxContactsReported(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_max_contacts_reported_(body)
}

fn physicsserver2dextension_gd_body_set_contacts_reported_depth_threshold[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetContactsReportedDepthThreshold(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	threshold := unsafe{&f64(args[1])}
	v_inst.body_set_contacts_reported_depth_threshold_(body, threshold)
}

fn physicsserver2dextension_gd_body_get_contacts_reported_depth_threshold[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetContactsReportedDepthThreshold(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.body_get_contacts_reported_depth_threshold_(body)
}

fn physicsserver2dextension_gd_body_set_omit_force_integration[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetOmitForceIntegration(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	enable := unsafe{&bool(args[1])}
	v_inst.body_set_omit_force_integration_(body, enable)
}

fn physicsserver2dextension_gd_body_is_omitting_force_integration[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyIsOmittingForceIntegration(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.body_is_omitting_force_integration_(body)
}

fn physicsserver2dextension_gd_body_set_state_sync_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetStateSyncCallback(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	callable := unsafe{&Callable(args[1])}
	v_inst.body_set_state_sync_callback_(body, callable)
}

fn physicsserver2dextension_gd_body_set_force_integration_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetForceIntegrationCallback(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	callable := unsafe{&Callable(args[1])}
	userdata := unsafe{&Variant(args[2])}
	v_inst.body_set_force_integration_callback_(body, callable, userdata)
}

fn physicsserver2dextension_gd_body_collide_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyCollideShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	body_shape := unsafe{&i64(args[1])}
	shape := unsafe{&RID(args[2])}
	shape_xform := unsafe{&Transform2D(args[3])}
	motion := unsafe{&Vector2(args[4])}
	results := unsafe{&voidptr(args[5])}
	result_max := unsafe{&i64(args[6])}
	result_count := unsafe{&&i32(args[7])}
	*(&bool(ret)) := v_inst.body_collide_shape_(body, body_shape, shape, shape_xform, motion, results, result_max, result_count)
}

fn physicsserver2dextension_gd_body_set_pickable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodySetPickable(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	pickable := unsafe{&bool(args[1])}
	v_inst.body_set_pickable_(body, pickable)
}

fn physicsserver2dextension_gd_body_get_direct_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyGetDirectState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&PhysicsDirectBodyState2D(ret)) := v_inst.body_get_direct_state_(body)
}

fn physicsserver2dextension_gd_body_test_motion[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionBodyTestMotion(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	from := unsafe{&Transform2D(args[1])}
	motion := unsafe{&Vector2(args[2])}
	margin := unsafe{&f64(args[3])}
	collide_separation_ray := unsafe{&bool(args[4])}
	recovery_as_collision := unsafe{&bool(args[5])}
	gd_result := unsafe{&&PhysicsServer2DExtensionMotionResult(args[6])}
	*(&bool(ret)) := v_inst.body_test_motion_(body, from, motion, margin, collide_separation_ray, recovery_as_collision, gd_result)
}

fn physicsserver2dextension_gd_joint_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.joint_create_()
}

fn physicsserver2dextension_gd_joint_clear[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointClear(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	v_inst.joint_clear_(joint)
}

fn physicsserver2dextension_gd_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DJointParam(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.joint_set_param_(joint, param, value)
}

fn physicsserver2dextension_gd_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DJointParam(args[1])}
	*(&f64(ret)) := v_inst.joint_get_param_(joint, param)
}

fn physicsserver2dextension_gd_joint_disable_collisions_between_bodies[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointDisableCollisionsBetweenBodies(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	disable := unsafe{&bool(args[1])}
	v_inst.joint_disable_collisions_between_bodies_(joint, disable)
}

fn physicsserver2dextension_gd_joint_is_disabled_collisions_between_bodies[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointIsDisabledCollisionsBetweenBodies(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.joint_is_disabled_collisions_between_bodies_(joint)
}

fn physicsserver2dextension_gd_joint_make_pin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointMakePin(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	anchor := unsafe{&Vector2(args[1])}
	body_a := unsafe{&RID(args[2])}
	body_b := unsafe{&RID(args[3])}
	v_inst.joint_make_pin_(joint, anchor, body_a, body_b)
}

fn physicsserver2dextension_gd_joint_make_groove[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointMakeGroove(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	a_groove1 := unsafe{&Vector2(args[1])}
	a_groove2 := unsafe{&Vector2(args[2])}
	b_anchor := unsafe{&Vector2(args[3])}
	body_a := unsafe{&RID(args[4])}
	body_b := unsafe{&RID(args[5])}
	v_inst.joint_make_groove_(joint, a_groove1, a_groove2, b_anchor, body_a, body_b)
}

fn physicsserver2dextension_gd_joint_make_damped_spring[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointMakeDampedSpring(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	anchor_a := unsafe{&Vector2(args[1])}
	anchor_b := unsafe{&Vector2(args[2])}
	body_a := unsafe{&RID(args[3])}
	body_b := unsafe{&RID(args[4])}
	v_inst.joint_make_damped_spring_(joint, anchor_a, anchor_b, body_a, body_b)
}

fn physicsserver2dextension_gd_pin_joint_set_flag[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionPinJointSetFlag(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	flag := unsafe{&PhysicsServer2DPinJointFlag(args[1])}
	enabled := unsafe{&bool(args[2])}
	v_inst.pin_joint_set_flag_(joint, flag, enabled)
}

fn physicsserver2dextension_gd_pin_joint_get_flag[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionPinJointGetFlag(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	flag := unsafe{&PhysicsServer2DPinJointFlag(args[1])}
	*(&bool(ret)) := v_inst.pin_joint_get_flag_(joint, flag)
}

fn physicsserver2dextension_gd_pin_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionPinJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DPinJointParam(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.pin_joint_set_param_(joint, param, value)
}

fn physicsserver2dextension_gd_pin_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionPinJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DPinJointParam(args[1])}
	*(&f64(ret)) := v_inst.pin_joint_get_param_(joint, param)
}

fn physicsserver2dextension_gd_damped_spring_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionDampedSpringJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DDampedSpringParam(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.damped_spring_joint_set_param_(joint, param, value)
}

fn physicsserver2dextension_gd_damped_spring_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionDampedSpringJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer2DDampedSpringParam(args[1])}
	*(&f64(ret)) := v_inst.damped_spring_joint_get_param_(joint, param)
}

fn physicsserver2dextension_gd_joint_get_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionJointGetType(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	*(&PhysicsServer2DJointType(ret)) := v_inst.joint_get_type_(joint)
}

fn physicsserver2dextension_gd_free_rid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionFreeRid(unsafe{&T(voidptr(inst))})
	rid := unsafe{&RID(args[0])}
	v_inst.free_rid_(rid)
}

fn physicsserver2dextension_gd_set_active[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSetActive(unsafe{&T(voidptr(inst))})
	active := unsafe{&bool(args[0])}
	v_inst.set_active_(active)
}

fn physicsserver2dextension_gd_init[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionInit(unsafe{&T(voidptr(inst))})
	v_inst.init_()
}

fn physicsserver2dextension_gd_step[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionStep(unsafe{&T(voidptr(inst))})
	step := unsafe{&f64(args[0])}
	v_inst.step_(step)
}

fn physicsserver2dextension_gd_sync[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionSync(unsafe{&T(voidptr(inst))})
	v_inst.sync_()
}

fn physicsserver2dextension_gd_flush_queries[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionFlushQueries(unsafe{&T(voidptr(inst))})
	v_inst.flush_queries_()
}

fn physicsserver2dextension_gd_end_sync[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionEndSync(unsafe{&T(voidptr(inst))})
	v_inst.end_sync_()
}

fn physicsserver2dextension_gd_finish[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionFinish(unsafe{&T(voidptr(inst))})
	v_inst.finish_()
}

fn physicsserver2dextension_gd_is_flushing_queries[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionIsFlushingQueries(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_flushing_queries_()
}

fn physicsserver2dextension_gd_get_process_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer2DExtensionGetProcessInfo(unsafe{&T(voidptr(inst))})
	process_info := unsafe{&PhysicsServer2DProcessInfo(args[0])}
	*(&i64(ret)) := v_inst.get_process_info_(process_info)
}

fn physicsserver3dextension_gd_world_boundary_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionWorldBoundaryShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.world_boundary_shape_create_()
}

fn physicsserver3dextension_gd_separation_ray_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSeparationRayShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.separation_ray_shape_create_()
}

fn physicsserver3dextension_gd_sphere_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSphereShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.sphere_shape_create_()
}

fn physicsserver3dextension_gd_box_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBoxShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.box_shape_create_()
}

fn physicsserver3dextension_gd_capsule_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionCapsuleShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.capsule_shape_create_()
}

fn physicsserver3dextension_gd_cylinder_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionCylinderShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.cylinder_shape_create_()
}

fn physicsserver3dextension_gd_convex_polygon_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionConvexPolygonShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.convex_polygon_shape_create_()
}

fn physicsserver3dextension_gd_concave_polygon_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionConcavePolygonShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.concave_polygon_shape_create_()
}

fn physicsserver3dextension_gd_heightmap_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionHeightmapShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.heightmap_shape_create_()
}

fn physicsserver3dextension_gd_custom_shape_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionCustomShapeCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.custom_shape_create_()
}

fn physicsserver3dextension_gd_shape_set_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionShapeSetData(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	data := unsafe{&Variant(args[1])}
	v_inst.shape_set_data_(shape, data)
}

fn physicsserver3dextension_gd_shape_set_custom_solver_bias[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionShapeSetCustomSolverBias(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	bias := unsafe{&f64(args[1])}
	v_inst.shape_set_custom_solver_bias_(shape, bias)
}

fn physicsserver3dextension_gd_shape_set_margin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionShapeSetMargin(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	margin := unsafe{&f64(args[1])}
	v_inst.shape_set_margin_(shape, margin)
}

fn physicsserver3dextension_gd_shape_get_margin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionShapeGetMargin(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shape_get_margin_(shape)
}

fn physicsserver3dextension_gd_shape_get_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionShapeGetType(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	*(&PhysicsServer3DShapeType(ret)) := v_inst.shape_get_type_(shape)
}

fn physicsserver3dextension_gd_shape_get_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionShapeGetData(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	*(&Variant(ret)) := v_inst.shape_get_data_(shape)
}

fn physicsserver3dextension_gd_shape_get_custom_solver_bias[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionShapeGetCustomSolverBias(unsafe{&T(voidptr(inst))})
	shape := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shape_get_custom_solver_bias_(shape)
}

fn physicsserver3dextension_gd_space_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.space_create_()
}

fn physicsserver3dextension_gd_space_set_active[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceSetActive(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	active := unsafe{&bool(args[1])}
	v_inst.space_set_active_(space, active)
}

fn physicsserver3dextension_gd_space_is_active[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceIsActive(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.space_is_active_(space)
}

fn physicsserver3dextension_gd_space_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceSetParam(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DSpaceParameter(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.space_set_param_(space, param, value)
}

fn physicsserver3dextension_gd_space_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceGetParam(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DSpaceParameter(args[1])}
	*(&f64(ret)) := v_inst.space_get_param_(space, param)
}

fn physicsserver3dextension_gd_space_get_direct_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceGetDirectState(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&PhysicsDirectSpaceState3D(ret)) := v_inst.space_get_direct_state_(space)
}

fn physicsserver3dextension_gd_space_set_debug_contacts[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceSetDebugContacts(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	max_contacts := unsafe{&i64(args[1])}
	v_inst.space_set_debug_contacts_(space, max_contacts)
}

fn physicsserver3dextension_gd_space_get_contacts[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceGetContacts(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&PackedVector3Array(ret)) := v_inst.space_get_contacts_(space)
}

fn physicsserver3dextension_gd_space_get_contact_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSpaceGetContactCount(unsafe{&T(voidptr(inst))})
	space := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.space_get_contact_count_(space)
}

fn physicsserver3dextension_gd_area_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.area_create_()
}

fn physicsserver3dextension_gd_area_set_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetSpace(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	space := unsafe{&RID(args[1])}
	v_inst.area_set_space_(area, space)
}

fn physicsserver3dextension_gd_area_get_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetSpace(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&RID(ret)) := v_inst.area_get_space_(area)
}

fn physicsserver3dextension_gd_area_add_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaAddShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape := unsafe{&RID(args[1])}
	transform := unsafe{&Transform3D(args[2])}
	disabled := unsafe{&bool(args[3])}
	v_inst.area_add_shape_(area, shape, transform, disabled)
}

fn physicsserver3dextension_gd_area_set_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	shape := unsafe{&RID(args[2])}
	v_inst.area_set_shape_(area, shape_idx, shape)
}

fn physicsserver3dextension_gd_area_set_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetShapeTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	transform := unsafe{&Transform3D(args[2])}
	v_inst.area_set_shape_transform_(area, shape_idx, transform)
}

fn physicsserver3dextension_gd_area_set_shape_disabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetShapeDisabled(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	disabled := unsafe{&bool(args[2])}
	v_inst.area_set_shape_disabled_(area, shape_idx, disabled)
}

fn physicsserver3dextension_gd_area_get_shape_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetShapeCount(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_shape_count_(area)
}

fn physicsserver3dextension_gd_area_get_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&RID(ret)) := v_inst.area_get_shape_(area, shape_idx)
}

fn physicsserver3dextension_gd_area_get_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetShapeTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&Transform3D(ret)) := v_inst.area_get_shape_transform_(area, shape_idx)
}

fn physicsserver3dextension_gd_area_remove_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaRemoveShape(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	v_inst.area_remove_shape_(area, shape_idx)
}

fn physicsserver3dextension_gd_area_clear_shapes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaClearShapes(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	v_inst.area_clear_shapes_(area)
}

fn physicsserver3dextension_gd_area_attach_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaAttachObjectInstanceId(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	id := unsafe{&i64(args[1])}
	v_inst.area_attach_object_instance_id_(area, id)
}

fn physicsserver3dextension_gd_area_get_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetObjectInstanceId(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_object_instance_id_(area)
}

fn physicsserver3dextension_gd_area_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetParam(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DAreaParameter(args[1])}
	value := unsafe{&Variant(args[2])}
	v_inst.area_set_param_(area, param, value)
}

fn physicsserver3dextension_gd_area_set_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	transform := unsafe{&Transform3D(args[1])}
	v_inst.area_set_transform_(area, transform)
}

fn physicsserver3dextension_gd_area_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetParam(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DAreaParameter(args[1])}
	*(&Variant(ret)) := v_inst.area_get_param_(area, param)
}

fn physicsserver3dextension_gd_area_get_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetTransform(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&Transform3D(ret)) := v_inst.area_get_transform_(area)
}

fn physicsserver3dextension_gd_area_set_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetCollisionLayer(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	layer := unsafe{&i64(args[1])}
	v_inst.area_set_collision_layer_(area, layer)
}

fn physicsserver3dextension_gd_area_get_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetCollisionLayer(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_collision_layer_(area)
}

fn physicsserver3dextension_gd_area_set_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetCollisionMask(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	mask := unsafe{&i64(args[1])}
	v_inst.area_set_collision_mask_(area, mask)
}

fn physicsserver3dextension_gd_area_get_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaGetCollisionMask(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.area_get_collision_mask_(area)
}

fn physicsserver3dextension_gd_area_set_monitorable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetMonitorable(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	monitorable := unsafe{&bool(args[1])}
	v_inst.area_set_monitorable_(area, monitorable)
}

fn physicsserver3dextension_gd_area_set_ray_pickable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetRayPickable(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	enable := unsafe{&bool(args[1])}
	v_inst.area_set_ray_pickable_(area, enable)
}

fn physicsserver3dextension_gd_area_set_monitor_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetMonitorCallback(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	callback := unsafe{&Callable(args[1])}
	v_inst.area_set_monitor_callback_(area, callback)
}

fn physicsserver3dextension_gd_area_set_area_monitor_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionAreaSetAreaMonitorCallback(unsafe{&T(voidptr(inst))})
	area := unsafe{&RID(args[0])}
	callback := unsafe{&Callable(args[1])}
	v_inst.area_set_area_monitor_callback_(area, callback)
}

fn physicsserver3dextension_gd_body_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.body_create_()
}

fn physicsserver3dextension_gd_body_set_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetSpace(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	space := unsafe{&RID(args[1])}
	v_inst.body_set_space_(body, space)
}

fn physicsserver3dextension_gd_body_get_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetSpace(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&RID(ret)) := v_inst.body_get_space_(body)
}

fn physicsserver3dextension_gd_body_set_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetMode(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	mode := unsafe{&PhysicsServer3DBodyMode(args[1])}
	v_inst.body_set_mode_(body, mode)
}

fn physicsserver3dextension_gd_body_get_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetMode(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&PhysicsServer3DBodyMode(ret)) := v_inst.body_get_mode_(body)
}

fn physicsserver3dextension_gd_body_add_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyAddShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape := unsafe{&RID(args[1])}
	transform := unsafe{&Transform3D(args[2])}
	disabled := unsafe{&bool(args[3])}
	v_inst.body_add_shape_(body, shape, transform, disabled)
}

fn physicsserver3dextension_gd_body_set_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	shape := unsafe{&RID(args[2])}
	v_inst.body_set_shape_(body, shape_idx, shape)
}

fn physicsserver3dextension_gd_body_set_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetShapeTransform(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	transform := unsafe{&Transform3D(args[2])}
	v_inst.body_set_shape_transform_(body, shape_idx, transform)
}

fn physicsserver3dextension_gd_body_set_shape_disabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetShapeDisabled(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	disabled := unsafe{&bool(args[2])}
	v_inst.body_set_shape_disabled_(body, shape_idx, disabled)
}

fn physicsserver3dextension_gd_body_get_shape_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetShapeCount(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_shape_count_(body)
}

fn physicsserver3dextension_gd_body_get_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&RID(ret)) := v_inst.body_get_shape_(body, shape_idx)
}

fn physicsserver3dextension_gd_body_get_shape_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetShapeTransform(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	*(&Transform3D(ret)) := v_inst.body_get_shape_transform_(body, shape_idx)
}

fn physicsserver3dextension_gd_body_remove_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyRemoveShape(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	shape_idx := unsafe{&i64(args[1])}
	v_inst.body_remove_shape_(body, shape_idx)
}

fn physicsserver3dextension_gd_body_clear_shapes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyClearShapes(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	v_inst.body_clear_shapes_(body)
}

fn physicsserver3dextension_gd_body_attach_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyAttachObjectInstanceId(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	id := unsafe{&i64(args[1])}
	v_inst.body_attach_object_instance_id_(body, id)
}

fn physicsserver3dextension_gd_body_get_object_instance_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetObjectInstanceId(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_object_instance_id_(body)
}

fn physicsserver3dextension_gd_body_set_enable_continuous_collision_detection[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetEnableContinuousCollisionDetection(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	enable := unsafe{&bool(args[1])}
	v_inst.body_set_enable_continuous_collision_detection_(body, enable)
}

fn physicsserver3dextension_gd_body_is_continuous_collision_detection_enabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyIsContinuousCollisionDetectionEnabled(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.body_is_continuous_collision_detection_enabled_(body)
}

fn physicsserver3dextension_gd_body_set_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetCollisionLayer(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	layer := unsafe{&i64(args[1])}
	v_inst.body_set_collision_layer_(body, layer)
}

fn physicsserver3dextension_gd_body_get_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetCollisionLayer(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_collision_layer_(body)
}

fn physicsserver3dextension_gd_body_set_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetCollisionMask(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	mask := unsafe{&i64(args[1])}
	v_inst.body_set_collision_mask_(body, mask)
}

fn physicsserver3dextension_gd_body_get_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetCollisionMask(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_collision_mask_(body)
}

fn physicsserver3dextension_gd_body_set_collision_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetCollisionPriority(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	priority := unsafe{&f64(args[1])}
	v_inst.body_set_collision_priority_(body, priority)
}

fn physicsserver3dextension_gd_body_get_collision_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetCollisionPriority(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.body_get_collision_priority_(body)
}

fn physicsserver3dextension_gd_body_set_user_flags[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetUserFlags(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	flags := unsafe{&i64(args[1])}
	v_inst.body_set_user_flags_(body, flags)
}

fn physicsserver3dextension_gd_body_get_user_flags[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetUserFlags(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_user_flags_(body)
}

fn physicsserver3dextension_gd_body_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetParam(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DBodyParameter(args[1])}
	value := unsafe{&Variant(args[2])}
	v_inst.body_set_param_(body, param, value)
}

fn physicsserver3dextension_gd_body_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetParam(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DBodyParameter(args[1])}
	*(&Variant(ret)) := v_inst.body_get_param_(body, param)
}

fn physicsserver3dextension_gd_body_reset_mass_properties[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyResetMassProperties(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	v_inst.body_reset_mass_properties_(body)
}

fn physicsserver3dextension_gd_body_set_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	state := unsafe{&PhysicsServer3DBodyState(args[1])}
	value := unsafe{&Variant(args[2])}
	v_inst.body_set_state_(body, state, value)
}

fn physicsserver3dextension_gd_body_get_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	state := unsafe{&PhysicsServer3DBodyState(args[1])}
	*(&Variant(ret)) := v_inst.body_get_state_(body, state)
}

fn physicsserver3dextension_gd_body_apply_central_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyApplyCentralImpulse(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	impulse := unsafe{&Vector3(args[1])}
	v_inst.body_apply_central_impulse_(body, impulse)
}

fn physicsserver3dextension_gd_body_apply_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyApplyImpulse(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	impulse := unsafe{&Vector3(args[1])}
	position := unsafe{&Vector3(args[2])}
	v_inst.body_apply_impulse_(body, impulse, position)
}

fn physicsserver3dextension_gd_body_apply_torque_impulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyApplyTorqueImpulse(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	impulse := unsafe{&Vector3(args[1])}
	v_inst.body_apply_torque_impulse_(body, impulse)
}

fn physicsserver3dextension_gd_body_apply_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyApplyCentralForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector3(args[1])}
	v_inst.body_apply_central_force_(body, force)
}

fn physicsserver3dextension_gd_body_apply_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyApplyForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector3(args[1])}
	position := unsafe{&Vector3(args[2])}
	v_inst.body_apply_force_(body, force, position)
}

fn physicsserver3dextension_gd_body_apply_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyApplyTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	torque := unsafe{&Vector3(args[1])}
	v_inst.body_apply_torque_(body, torque)
}

fn physicsserver3dextension_gd_body_add_constant_central_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyAddConstantCentralForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector3(args[1])}
	v_inst.body_add_constant_central_force_(body, force)
}

fn physicsserver3dextension_gd_body_add_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyAddConstantForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector3(args[1])}
	position := unsafe{&Vector3(args[2])}
	v_inst.body_add_constant_force_(body, force, position)
}

fn physicsserver3dextension_gd_body_add_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyAddConstantTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	torque := unsafe{&Vector3(args[1])}
	v_inst.body_add_constant_torque_(body, torque)
}

fn physicsserver3dextension_gd_body_set_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetConstantForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	force := unsafe{&Vector3(args[1])}
	v_inst.body_set_constant_force_(body, force)
}

fn physicsserver3dextension_gd_body_get_constant_force[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetConstantForce(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&Vector3(ret)) := v_inst.body_get_constant_force_(body)
}

fn physicsserver3dextension_gd_body_set_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetConstantTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	torque := unsafe{&Vector3(args[1])}
	v_inst.body_set_constant_torque_(body, torque)
}

fn physicsserver3dextension_gd_body_get_constant_torque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetConstantTorque(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&Vector3(ret)) := v_inst.body_get_constant_torque_(body)
}

fn physicsserver3dextension_gd_body_set_axis_velocity[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetAxisVelocity(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	axis_velocity := unsafe{&Vector3(args[1])}
	v_inst.body_set_axis_velocity_(body, axis_velocity)
}

fn physicsserver3dextension_gd_body_set_axis_lock[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetAxisLock(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	axis := unsafe{&PhysicsServer3DBodyAxis(args[1])}
	gd_lock := unsafe{&bool(args[2])}
	v_inst.body_set_axis_lock_(body, axis, gd_lock)
}

fn physicsserver3dextension_gd_body_is_axis_locked[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyIsAxisLocked(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	axis := unsafe{&PhysicsServer3DBodyAxis(args[1])}
	*(&bool(ret)) := v_inst.body_is_axis_locked_(body, axis)
}

fn physicsserver3dextension_gd_body_add_collision_exception[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyAddCollisionException(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	excepted_body := unsafe{&RID(args[1])}
	v_inst.body_add_collision_exception_(body, excepted_body)
}

fn physicsserver3dextension_gd_body_remove_collision_exception[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyRemoveCollisionException(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	excepted_body := unsafe{&RID(args[1])}
	v_inst.body_remove_collision_exception_(body, excepted_body)
}

fn physicsserver3dextension_gd_body_get_collision_exceptions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetCollisionExceptions(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&Array(ret)) := v_inst.body_get_collision_exceptions_(body)
}

fn physicsserver3dextension_gd_body_set_max_contacts_reported[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetMaxContactsReported(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	amount := unsafe{&i64(args[1])}
	v_inst.body_set_max_contacts_reported_(body, amount)
}

fn physicsserver3dextension_gd_body_get_max_contacts_reported[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetMaxContactsReported(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.body_get_max_contacts_reported_(body)
}

fn physicsserver3dextension_gd_body_set_contacts_reported_depth_threshold[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetContactsReportedDepthThreshold(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	threshold := unsafe{&f64(args[1])}
	v_inst.body_set_contacts_reported_depth_threshold_(body, threshold)
}

fn physicsserver3dextension_gd_body_get_contacts_reported_depth_threshold[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetContactsReportedDepthThreshold(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.body_get_contacts_reported_depth_threshold_(body)
}

fn physicsserver3dextension_gd_body_set_omit_force_integration[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetOmitForceIntegration(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	enable := unsafe{&bool(args[1])}
	v_inst.body_set_omit_force_integration_(body, enable)
}

fn physicsserver3dextension_gd_body_is_omitting_force_integration[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyIsOmittingForceIntegration(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.body_is_omitting_force_integration_(body)
}

fn physicsserver3dextension_gd_body_set_state_sync_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetStateSyncCallback(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	callable := unsafe{&Callable(args[1])}
	v_inst.body_set_state_sync_callback_(body, callable)
}

fn physicsserver3dextension_gd_body_set_force_integration_callback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetForceIntegrationCallback(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	callable := unsafe{&Callable(args[1])}
	userdata := unsafe{&Variant(args[2])}
	v_inst.body_set_force_integration_callback_(body, callable, userdata)
}

fn physicsserver3dextension_gd_body_set_ray_pickable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodySetRayPickable(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	enable := unsafe{&bool(args[1])}
	v_inst.body_set_ray_pickable_(body, enable)
}

fn physicsserver3dextension_gd_body_test_motion[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyTestMotion(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	from := unsafe{&Transform3D(args[1])}
	motion := unsafe{&Vector3(args[2])}
	margin := unsafe{&f64(args[3])}
	max_collisions := unsafe{&i64(args[4])}
	collide_separation_ray := unsafe{&bool(args[5])}
	recovery_as_collision := unsafe{&bool(args[6])}
	gd_result := unsafe{&&PhysicsServer3DExtensionMotionResult(args[7])}
	*(&bool(ret)) := v_inst.body_test_motion_(body, from, motion, margin, max_collisions, collide_separation_ray, recovery_as_collision, gd_result)
}

fn physicsserver3dextension_gd_body_get_direct_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionBodyGetDirectState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&PhysicsDirectBodyState3D(ret)) := v_inst.body_get_direct_state_(body)
}

fn physicsserver3dextension_gd_soft_body_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.soft_body_create_()
}

fn physicsserver3dextension_gd_soft_body_update_rendering_server[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyUpdateRenderingServer(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	rendering_server_handler := unsafe{&PhysicsServer3DRenderingServerHandler(args[1])}
	v_inst.soft_body_update_rendering_server_(body, rendering_server_handler)
}

fn physicsserver3dextension_gd_soft_body_set_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetSpace(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	space := unsafe{&RID(args[1])}
	v_inst.soft_body_set_space_(body, space)
}

fn physicsserver3dextension_gd_soft_body_get_space[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetSpace(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&RID(ret)) := v_inst.soft_body_get_space_(body)
}

fn physicsserver3dextension_gd_soft_body_set_ray_pickable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetRayPickable(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	enable := unsafe{&bool(args[1])}
	v_inst.soft_body_set_ray_pickable_(body, enable)
}

fn physicsserver3dextension_gd_soft_body_set_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetCollisionLayer(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	layer := unsafe{&i64(args[1])}
	v_inst.soft_body_set_collision_layer_(body, layer)
}

fn physicsserver3dextension_gd_soft_body_get_collision_layer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetCollisionLayer(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.soft_body_get_collision_layer_(body)
}

fn physicsserver3dextension_gd_soft_body_set_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetCollisionMask(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	mask := unsafe{&i64(args[1])}
	v_inst.soft_body_set_collision_mask_(body, mask)
}

fn physicsserver3dextension_gd_soft_body_get_collision_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetCollisionMask(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.soft_body_get_collision_mask_(body)
}

fn physicsserver3dextension_gd_soft_body_add_collision_exception[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyAddCollisionException(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	body_b := unsafe{&RID(args[1])}
	v_inst.soft_body_add_collision_exception_(body, body_b)
}

fn physicsserver3dextension_gd_soft_body_remove_collision_exception[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyRemoveCollisionException(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	body_b := unsafe{&RID(args[1])}
	v_inst.soft_body_remove_collision_exception_(body, body_b)
}

fn physicsserver3dextension_gd_soft_body_get_collision_exceptions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetCollisionExceptions(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&Array(ret)) := v_inst.soft_body_get_collision_exceptions_(body)
}

fn physicsserver3dextension_gd_soft_body_set_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	state := unsafe{&PhysicsServer3DBodyState(args[1])}
	variant := unsafe{&Variant(args[2])}
	v_inst.soft_body_set_state_(body, state, variant)
}

fn physicsserver3dextension_gd_soft_body_get_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetState(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	state := unsafe{&PhysicsServer3DBodyState(args[1])}
	*(&Variant(ret)) := v_inst.soft_body_get_state_(body, state)
}

fn physicsserver3dextension_gd_soft_body_set_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetTransform(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	transform := unsafe{&Transform3D(args[1])}
	v_inst.soft_body_set_transform_(body, transform)
}

fn physicsserver3dextension_gd_soft_body_set_simulation_precision[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetSimulationPrecision(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	simulation_precision := unsafe{&i64(args[1])}
	v_inst.soft_body_set_simulation_precision_(body, simulation_precision)
}

fn physicsserver3dextension_gd_soft_body_get_simulation_precision[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetSimulationPrecision(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.soft_body_get_simulation_precision_(body)
}

fn physicsserver3dextension_gd_soft_body_set_total_mass[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetTotalMass(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	total_mass := unsafe{&f64(args[1])}
	v_inst.soft_body_set_total_mass_(body, total_mass)
}

fn physicsserver3dextension_gd_soft_body_get_total_mass[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetTotalMass(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.soft_body_get_total_mass_(body)
}

fn physicsserver3dextension_gd_soft_body_set_linear_stiffness[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetLinearStiffness(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	linear_stiffness := unsafe{&f64(args[1])}
	v_inst.soft_body_set_linear_stiffness_(body, linear_stiffness)
}

fn physicsserver3dextension_gd_soft_body_get_linear_stiffness[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetLinearStiffness(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.soft_body_get_linear_stiffness_(body)
}

fn physicsserver3dextension_gd_soft_body_set_pressure_coefficient[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetPressureCoefficient(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	pressure_coefficient := unsafe{&f64(args[1])}
	v_inst.soft_body_set_pressure_coefficient_(body, pressure_coefficient)
}

fn physicsserver3dextension_gd_soft_body_get_pressure_coefficient[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetPressureCoefficient(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.soft_body_get_pressure_coefficient_(body)
}

fn physicsserver3dextension_gd_soft_body_set_damping_coefficient[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetDampingCoefficient(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	damping_coefficient := unsafe{&f64(args[1])}
	v_inst.soft_body_set_damping_coefficient_(body, damping_coefficient)
}

fn physicsserver3dextension_gd_soft_body_get_damping_coefficient[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetDampingCoefficient(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.soft_body_get_damping_coefficient_(body)
}

fn physicsserver3dextension_gd_soft_body_set_drag_coefficient[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetDragCoefficient(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	drag_coefficient := unsafe{&f64(args[1])}
	v_inst.soft_body_set_drag_coefficient_(body, drag_coefficient)
}

fn physicsserver3dextension_gd_soft_body_get_drag_coefficient[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetDragCoefficient(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.soft_body_get_drag_coefficient_(body)
}

fn physicsserver3dextension_gd_soft_body_set_mesh[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodySetMesh(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	mesh := unsafe{&RID(args[1])}
	v_inst.soft_body_set_mesh_(body, mesh)
}

fn physicsserver3dextension_gd_soft_body_get_bounds[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetBounds(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	*(&AABB(ret)) := v_inst.soft_body_get_bounds_(body)
}

fn physicsserver3dextension_gd_soft_body_move_point[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyMovePoint(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	point_index := unsafe{&i64(args[1])}
	global_position := unsafe{&Vector3(args[2])}
	v_inst.soft_body_move_point_(body, point_index, global_position)
}

fn physicsserver3dextension_gd_soft_body_get_point_global_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyGetPointGlobalPosition(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	point_index := unsafe{&i64(args[1])}
	*(&Vector3(ret)) := v_inst.soft_body_get_point_global_position_(body, point_index)
}

fn physicsserver3dextension_gd_soft_body_remove_all_pinned_points[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyRemoveAllPinnedPoints(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	v_inst.soft_body_remove_all_pinned_points_(body)
}

fn physicsserver3dextension_gd_soft_body_pin_point[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyPinPoint(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	point_index := unsafe{&i64(args[1])}
	pin := unsafe{&bool(args[2])}
	v_inst.soft_body_pin_point_(body, point_index, pin)
}

fn physicsserver3dextension_gd_soft_body_is_point_pinned[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSoftBodyIsPointPinned(unsafe{&T(voidptr(inst))})
	body := unsafe{&RID(args[0])}
	point_index := unsafe{&i64(args[1])}
	*(&bool(ret)) := v_inst.soft_body_is_point_pinned_(body, point_index)
}

fn physicsserver3dextension_gd_joint_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointCreate(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.joint_create_()
}

fn physicsserver3dextension_gd_joint_clear[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointClear(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	v_inst.joint_clear_(joint)
}

fn physicsserver3dextension_gd_joint_make_pin[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointMakePin(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	body_a := unsafe{&RID(args[1])}
	local_a := unsafe{&Vector3(args[2])}
	body_b := unsafe{&RID(args[3])}
	local_b := unsafe{&Vector3(args[4])}
	v_inst.joint_make_pin_(joint, body_a, local_a, body_b, local_b)
}

fn physicsserver3dextension_gd_pin_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionPinJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DPinJointParam(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.pin_joint_set_param_(joint, param, value)
}

fn physicsserver3dextension_gd_pin_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionPinJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DPinJointParam(args[1])}
	*(&f64(ret)) := v_inst.pin_joint_get_param_(joint, param)
}

fn physicsserver3dextension_gd_pin_joint_set_local_a[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionPinJointSetLocalA(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	local_a := unsafe{&Vector3(args[1])}
	v_inst.pin_joint_set_local_a_(joint, local_a)
}

fn physicsserver3dextension_gd_pin_joint_get_local_a[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionPinJointGetLocalA(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	*(&Vector3(ret)) := v_inst.pin_joint_get_local_a_(joint)
}

fn physicsserver3dextension_gd_pin_joint_set_local_b[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionPinJointSetLocalB(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	local_b := unsafe{&Vector3(args[1])}
	v_inst.pin_joint_set_local_b_(joint, local_b)
}

fn physicsserver3dextension_gd_pin_joint_get_local_b[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionPinJointGetLocalB(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	*(&Vector3(ret)) := v_inst.pin_joint_get_local_b_(joint)
}

fn physicsserver3dextension_gd_joint_make_hinge[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointMakeHinge(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	body_a := unsafe{&RID(args[1])}
	hinge_a := unsafe{&Transform3D(args[2])}
	body_b := unsafe{&RID(args[3])}
	hinge_b := unsafe{&Transform3D(args[4])}
	v_inst.joint_make_hinge_(joint, body_a, hinge_a, body_b, hinge_b)
}

fn physicsserver3dextension_gd_joint_make_hinge_simple[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointMakeHingeSimple(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	body_a := unsafe{&RID(args[1])}
	pivot_a := unsafe{&Vector3(args[2])}
	axis_a := unsafe{&Vector3(args[3])}
	body_b := unsafe{&RID(args[4])}
	pivot_b := unsafe{&Vector3(args[5])}
	axis_b := unsafe{&Vector3(args[6])}
	v_inst.joint_make_hinge_simple_(joint, body_a, pivot_a, axis_a, body_b, pivot_b, axis_b)
}

fn physicsserver3dextension_gd_hinge_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionHingeJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DHingeJointParam(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.hinge_joint_set_param_(joint, param, value)
}

fn physicsserver3dextension_gd_hinge_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionHingeJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DHingeJointParam(args[1])}
	*(&f64(ret)) := v_inst.hinge_joint_get_param_(joint, param)
}

fn physicsserver3dextension_gd_hinge_joint_set_flag[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionHingeJointSetFlag(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	flag := unsafe{&PhysicsServer3DHingeJointFlag(args[1])}
	enabled := unsafe{&bool(args[2])}
	v_inst.hinge_joint_set_flag_(joint, flag, enabled)
}

fn physicsserver3dextension_gd_hinge_joint_get_flag[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionHingeJointGetFlag(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	flag := unsafe{&PhysicsServer3DHingeJointFlag(args[1])}
	*(&bool(ret)) := v_inst.hinge_joint_get_flag_(joint, flag)
}

fn physicsserver3dextension_gd_joint_make_slider[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointMakeSlider(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	body_a := unsafe{&RID(args[1])}
	local_ref_a := unsafe{&Transform3D(args[2])}
	body_b := unsafe{&RID(args[3])}
	local_ref_b := unsafe{&Transform3D(args[4])}
	v_inst.joint_make_slider_(joint, body_a, local_ref_a, body_b, local_ref_b)
}

fn physicsserver3dextension_gd_slider_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSliderJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DSliderJointParam(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.slider_joint_set_param_(joint, param, value)
}

fn physicsserver3dextension_gd_slider_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSliderJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DSliderJointParam(args[1])}
	*(&f64(ret)) := v_inst.slider_joint_get_param_(joint, param)
}

fn physicsserver3dextension_gd_joint_make_cone_twist[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointMakeConeTwist(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	body_a := unsafe{&RID(args[1])}
	local_ref_a := unsafe{&Transform3D(args[2])}
	body_b := unsafe{&RID(args[3])}
	local_ref_b := unsafe{&Transform3D(args[4])}
	v_inst.joint_make_cone_twist_(joint, body_a, local_ref_a, body_b, local_ref_b)
}

fn physicsserver3dextension_gd_cone_twist_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionConeTwistJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DConeTwistJointParam(args[1])}
	value := unsafe{&f64(args[2])}
	v_inst.cone_twist_joint_set_param_(joint, param, value)
}

fn physicsserver3dextension_gd_cone_twist_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionConeTwistJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	param := unsafe{&PhysicsServer3DConeTwistJointParam(args[1])}
	*(&f64(ret)) := v_inst.cone_twist_joint_get_param_(joint, param)
}

fn physicsserver3dextension_gd_joint_make_generic_6dof[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointMakeGeneric6dof(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	body_a := unsafe{&RID(args[1])}
	local_ref_a := unsafe{&Transform3D(args[2])}
	body_b := unsafe{&RID(args[3])}
	local_ref_b := unsafe{&Transform3D(args[4])}
	v_inst.joint_make_generic_6dof_(joint, body_a, local_ref_a, body_b, local_ref_b)
}

fn physicsserver3dextension_gd_generic_6dof_joint_set_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionGeneric6dofJointSetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	axis := unsafe{&Vector3Axis(args[1])}
	param := unsafe{&PhysicsServer3DG6DOFJointAxisParam(args[2])}
	value := unsafe{&f64(args[3])}
	v_inst.generic_6dof_joint_set_param_(joint, axis, param, value)
}

fn physicsserver3dextension_gd_generic_6dof_joint_get_param[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionGeneric6dofJointGetParam(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	axis := unsafe{&Vector3Axis(args[1])}
	param := unsafe{&PhysicsServer3DG6DOFJointAxisParam(args[2])}
	*(&f64(ret)) := v_inst.generic_6dof_joint_get_param_(joint, axis, param)
}

fn physicsserver3dextension_gd_generic_6dof_joint_set_flag[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionGeneric6dofJointSetFlag(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	axis := unsafe{&Vector3Axis(args[1])}
	flag := unsafe{&PhysicsServer3DG6DOFJointAxisFlag(args[2])}
	enable := unsafe{&bool(args[3])}
	v_inst.generic_6dof_joint_set_flag_(joint, axis, flag, enable)
}

fn physicsserver3dextension_gd_generic_6dof_joint_get_flag[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionGeneric6dofJointGetFlag(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	axis := unsafe{&Vector3Axis(args[1])}
	flag := unsafe{&PhysicsServer3DG6DOFJointAxisFlag(args[2])}
	*(&bool(ret)) := v_inst.generic_6dof_joint_get_flag_(joint, axis, flag)
}

fn physicsserver3dextension_gd_joint_get_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointGetType(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	*(&PhysicsServer3DJointType(ret)) := v_inst.joint_get_type_(joint)
}

fn physicsserver3dextension_gd_joint_set_solver_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointSetSolverPriority(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	priority := unsafe{&i64(args[1])}
	v_inst.joint_set_solver_priority_(joint, priority)
}

fn physicsserver3dextension_gd_joint_get_solver_priority[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointGetSolverPriority(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.joint_get_solver_priority_(joint)
}

fn physicsserver3dextension_gd_joint_disable_collisions_between_bodies[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointDisableCollisionsBetweenBodies(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	disable := unsafe{&bool(args[1])}
	v_inst.joint_disable_collisions_between_bodies_(joint, disable)
}

fn physicsserver3dextension_gd_joint_is_disabled_collisions_between_bodies[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionJointIsDisabledCollisionsBetweenBodies(unsafe{&T(voidptr(inst))})
	joint := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.joint_is_disabled_collisions_between_bodies_(joint)
}

fn physicsserver3dextension_gd_free_rid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionFreeRid(unsafe{&T(voidptr(inst))})
	rid := unsafe{&RID(args[0])}
	v_inst.free_rid_(rid)
}

fn physicsserver3dextension_gd_set_active[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSetActive(unsafe{&T(voidptr(inst))})
	active := unsafe{&bool(args[0])}
	v_inst.set_active_(active)
}

fn physicsserver3dextension_gd_init[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionInit(unsafe{&T(voidptr(inst))})
	v_inst.init_()
}

fn physicsserver3dextension_gd_step[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionStep(unsafe{&T(voidptr(inst))})
	step := unsafe{&f64(args[0])}
	v_inst.step_(step)
}

fn physicsserver3dextension_gd_sync[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionSync(unsafe{&T(voidptr(inst))})
	v_inst.sync_()
}

fn physicsserver3dextension_gd_flush_queries[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionFlushQueries(unsafe{&T(voidptr(inst))})
	v_inst.flush_queries_()
}

fn physicsserver3dextension_gd_end_sync[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionEndSync(unsafe{&T(voidptr(inst))})
	v_inst.end_sync_()
}

fn physicsserver3dextension_gd_finish[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionFinish(unsafe{&T(voidptr(inst))})
	v_inst.finish_()
}

fn physicsserver3dextension_gd_is_flushing_queries[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionIsFlushingQueries(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_flushing_queries_()
}

fn physicsserver3dextension_gd_get_process_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DExtensionGetProcessInfo(unsafe{&T(voidptr(inst))})
	process_info := unsafe{&PhysicsServer3DProcessInfo(args[0])}
	*(&i64(ret)) := v_inst.get_process_info_(process_info)
}

fn physicsserver3drenderingserverhandler_gd_set_vertex[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DRenderingServerHandlerSetVertex(unsafe{&T(voidptr(inst))})
	vertex_id := unsafe{&i64(args[0])}
	vertex := unsafe{&Vector3(args[1])}
	v_inst.set_vertex_(vertex_id, vertex)
}

fn physicsserver3drenderingserverhandler_gd_set_normal[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DRenderingServerHandlerSetNormal(unsafe{&T(voidptr(inst))})
	vertex_id := unsafe{&i64(args[0])}
	normal := unsafe{&Vector3(args[1])}
	v_inst.set_normal_(vertex_id, normal)
}

fn physicsserver3drenderingserverhandler_gd_set_aabb[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPhysicsServer3DRenderingServerHandlerSetAabb(unsafe{&T(voidptr(inst))})
	aabb := unsafe{&AABB(args[0])}
	v_inst.set_aabb_(aabb)
}

fn primitivemesh_gd_create_mesh_array[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IPrimitiveMeshCreateMeshArray(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.create_mesh_array_()
}

fn range_gd_value_changed[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRangeValueChanged(unsafe{&T(voidptr(inst))})
	new_value := unsafe{&f64(args[0])}
	v_inst.value_changed_(new_value)
}

fn renderdataextension_gd_get_render_scene_buffers[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderDataExtensionGetRenderSceneBuffers(unsafe{&T(voidptr(inst))})
	*(&RenderSceneBuffers(ret)) := v_inst.get_render_scene_buffers_()
}

fn renderdataextension_gd_get_render_scene_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderDataExtensionGetRenderSceneData(unsafe{&T(voidptr(inst))})
	*(&RenderSceneData(ret)) := v_inst.get_render_scene_data_()
}

fn renderdataextension_gd_get_environment[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderDataExtensionGetEnvironment(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_environment_()
}

fn renderdataextension_gd_get_camera_attributes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderDataExtensionGetCameraAttributes(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_camera_attributes_()
}

fn renderscenebuffersextension_gd_configure[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneBuffersExtensionConfigure(unsafe{&T(voidptr(inst))})
	config := unsafe{&RenderSceneBuffersConfiguration(args[0])}
	v_inst.configure_(config)
}

fn renderscenebuffersextension_gd_set_fsr_sharpness[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneBuffersExtensionSetFsrSharpness(unsafe{&T(voidptr(inst))})
	fsr_sharpness := unsafe{&f64(args[0])}
	v_inst.set_fsr_sharpness_(fsr_sharpness)
}

fn renderscenebuffersextension_gd_set_texture_mipmap_bias[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneBuffersExtensionSetTextureMipmapBias(unsafe{&T(voidptr(inst))})
	texture_mipmap_bias := unsafe{&f64(args[0])}
	v_inst.set_texture_mipmap_bias_(texture_mipmap_bias)
}

fn renderscenebuffersextension_gd_set_anisotropic_filtering_level[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneBuffersExtensionSetAnisotropicFilteringLevel(unsafe{&T(voidptr(inst))})
	anisotropic_filtering_level := unsafe{&i64(args[0])}
	v_inst.set_anisotropic_filtering_level_(anisotropic_filtering_level)
}

fn renderscenebuffersextension_gd_set_use_debanding[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneBuffersExtensionSetUseDebanding(unsafe{&T(voidptr(inst))})
	use_debanding := unsafe{&bool(args[0])}
	v_inst.set_use_debanding_(use_debanding)
}

fn renderscenedataextension_gd_get_cam_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneDataExtensionGetCamTransform(unsafe{&T(voidptr(inst))})
	*(&Transform3D(ret)) := v_inst.get_cam_transform_()
}

fn renderscenedataextension_gd_get_cam_projection[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneDataExtensionGetCamProjection(unsafe{&T(voidptr(inst))})
	*(&Projection(ret)) := v_inst.get_cam_projection_()
}

fn renderscenedataextension_gd_get_view_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneDataExtensionGetViewCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_view_count_()
}

fn renderscenedataextension_gd_get_view_eye_offset[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneDataExtensionGetViewEyeOffset(unsafe{&T(voidptr(inst))})
	view := unsafe{&i64(args[0])}
	*(&Vector3(ret)) := v_inst.get_view_eye_offset_(view)
}

fn renderscenedataextension_gd_get_view_projection[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneDataExtensionGetViewProjection(unsafe{&T(voidptr(inst))})
	view := unsafe{&i64(args[0])}
	*(&Projection(ret)) := v_inst.get_view_projection_(view)
}

fn renderscenedataextension_gd_get_uniform_buffer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRenderSceneDataExtensionGetUniformBuffer(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_uniform_buffer_()
}

fn resource_gd_setup_local_to_scene[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceSetupLocalToScene(unsafe{&T(voidptr(inst))})
	v_inst.setup_local_to_scene_()
}

fn resource_gd_get_rid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceGetRid(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_rid_()
}

fn resource_gd_reset_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceResetState(unsafe{&T(voidptr(inst))})
	v_inst.reset_state_()
}

fn resource_gd_set_path_cache[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceSetPathCache(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	v_inst.set_path_cache_(path)
}

fn resourceformatloader_gd_get_recognized_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderGetRecognizedExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_recognized_extensions_()
}

fn resourceformatloader_gd_recognize_path[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderRecognizePath(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	gd_type := unsafe{&StringName(args[1])}
	*(&bool(ret)) := v_inst.recognize_path_(path, gd_type)
}

fn resourceformatloader_gd_handles_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderHandlesType(unsafe{&T(voidptr(inst))})
	gd_type := unsafe{&StringName(args[0])}
	*(&bool(ret)) := v_inst.handles_type_(gd_type)
}

fn resourceformatloader_gd_get_resource_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderGetResourceType(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&String(ret)) := v_inst.get_resource_type_(path)
}

fn resourceformatloader_gd_get_resource_script_class[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderGetResourceScriptClass(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&String(ret)) := v_inst.get_resource_script_class_(path)
}

fn resourceformatloader_gd_get_resource_uid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderGetResourceUid(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&i64(ret)) := v_inst.get_resource_uid_(path)
}

fn resourceformatloader_gd_get_dependencies[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderGetDependencies(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	add_types := unsafe{&bool(args[1])}
	*(&PackedStringArray(ret)) := v_inst.get_dependencies_(path, add_types)
}

fn resourceformatloader_gd_rename_dependencies[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderRenameDependencies(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	renames := unsafe{&Dictionary(args[1])}
	*(&GDError(ret)) := v_inst.rename_dependencies_(path, renames)
}

fn resourceformatloader_gd_exists[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderExists(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.exists_(path)
}

fn resourceformatloader_gd_get_classes_used[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderGetClassesUsed(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&PackedStringArray(ret)) := v_inst.get_classes_used_(path)
}

fn resourceformatloader_gd_load[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatLoaderLoad(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	original_path := unsafe{&String(args[1])}
	use_sub_threads := unsafe{&bool(args[2])}
	cache_mode := unsafe{&i64(args[3])}
	*(&Variant(ret)) := v_inst.load_(path, original_path, use_sub_threads, cache_mode)
}

fn resourceformatsaver_gd_save[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatSaverSave(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	path := unsafe{&String(args[1])}
	flags := unsafe{&i64(args[2])}
	*(&GDError(ret)) := v_inst.save_(resource, path, flags)
}

fn resourceformatsaver_gd_set_uid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatSaverSetUid(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	uid := unsafe{&i64(args[1])}
	*(&GDError(ret)) := v_inst.set_uid_(path, uid)
}

fn resourceformatsaver_gd_recognize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatSaverRecognize(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	*(&bool(ret)) := v_inst.recognize_(resource)
}

fn resourceformatsaver_gd_get_recognized_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatSaverGetRecognizedExtensions(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	*(&PackedStringArray(ret)) := v_inst.get_recognized_extensions_(resource)
}

fn resourceformatsaver_gd_recognize_path[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IResourceFormatSaverRecognizePath(unsafe{&T(voidptr(inst))})
	resource := unsafe{&Resource(args[0])}
	path := unsafe{&String(args[1])}
	*(&bool(ret)) := v_inst.recognize_path_(resource, path)
}

fn richtexteffect_gd_process_custom_fx[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRichTextEffectProcessCustomFx(unsafe{&T(voidptr(inst))})
	char_fx := unsafe{&CharFXTransform(args[0])}
	*(&bool(ret)) := v_inst.process_custom_fx_(char_fx)
}

fn rigidbody2d_gd_integrate_forces[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRigidBody2DIntegrateForces(unsafe{&T(voidptr(inst))})
	state := unsafe{&PhysicsDirectBodyState2D(args[0])}
	v_inst.integrate_forces_(state)
}

fn rigidbody3d_gd_integrate_forces[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IRigidBody3DIntegrateForces(unsafe{&T(voidptr(inst))})
	state := unsafe{&PhysicsDirectBodyState3D(args[0])}
	v_inst.integrate_forces_(state)
}

fn scriptextension_gd_editor_can_reload_from_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionEditorCanReloadFromFile(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.editor_can_reload_from_file_()
}

fn scriptextension_gd_placeholder_erased[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionPlaceholderErased(unsafe{&T(voidptr(inst))})
	placeholder := unsafe{&voidptr(args[0])}
	v_inst.placeholder_erased_(placeholder)
}

fn scriptextension_gd_can_instantiate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionCanInstantiate(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_instantiate_()
}

fn scriptextension_gd_get_base_script[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetBaseScript(unsafe{&T(voidptr(inst))})
	*(&Script(ret)) := v_inst.get_base_script_()
}

fn scriptextension_gd_get_global_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetGlobalName(unsafe{&T(voidptr(inst))})
	*(&StringName(ret)) := v_inst.get_global_name_()
}

fn scriptextension_gd_inherits_script[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionInheritsScript(unsafe{&T(voidptr(inst))})
	script := unsafe{&Script(args[0])}
	*(&bool(ret)) := v_inst.inherits_script_(script)
}

fn scriptextension_gd_get_instance_base_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetInstanceBaseType(unsafe{&T(voidptr(inst))})
	*(&StringName(ret)) := v_inst.get_instance_base_type_()
}

fn scriptextension_gd_instance_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionInstanceCreate(unsafe{&T(voidptr(inst))})
	for_object := unsafe{&Object(args[0])}
	*(&voidptr(ret)) := v_inst.instance_create_(for_object)
}

fn scriptextension_gd_placeholder_instance_create[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionPlaceholderInstanceCreate(unsafe{&T(voidptr(inst))})
	for_object := unsafe{&Object(args[0])}
	*(&voidptr(ret)) := v_inst.placeholder_instance_create_(for_object)
}

fn scriptextension_gd_instance_has[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionInstanceHas(unsafe{&T(voidptr(inst))})
	object := unsafe{&Object(args[0])}
	*(&bool(ret)) := v_inst.instance_has_(object)
}

fn scriptextension_gd_has_source_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionHasSourceCode(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_source_code_()
}

fn scriptextension_gd_get_source_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetSourceCode(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_source_code_()
}

fn scriptextension_gd_set_source_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionSetSourceCode(unsafe{&T(voidptr(inst))})
	code := unsafe{&String(args[0])}
	v_inst.set_source_code_(code)
}

fn scriptextension_gd_reload[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionReload(unsafe{&T(voidptr(inst))})
	keep_state := unsafe{&bool(args[0])}
	*(&GDError(ret)) := v_inst.reload_(keep_state)
}

fn scriptextension_gd_get_doc_class_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetDocClassName(unsafe{&T(voidptr(inst))})
	*(&StringName(ret)) := v_inst.get_doc_class_name_()
}

fn scriptextension_gd_get_documentation[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetDocumentation(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_documentation_()
}

fn scriptextension_gd_get_class_icon_path[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetClassIconPath(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_class_icon_path_()
}

fn scriptextension_gd_has_method[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionHasMethod(unsafe{&T(voidptr(inst))})
	method := unsafe{&StringName(args[0])}
	*(&bool(ret)) := v_inst.has_method_(method)
}

fn scriptextension_gd_has_static_method[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionHasStaticMethod(unsafe{&T(voidptr(inst))})
	method := unsafe{&StringName(args[0])}
	*(&bool(ret)) := v_inst.has_static_method_(method)
}

fn scriptextension_gd_get_script_method_argument_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetScriptMethodArgumentCount(unsafe{&T(voidptr(inst))})
	method := unsafe{&StringName(args[0])}
	*(&Variant(ret)) := v_inst.get_script_method_argument_count_(method)
}

fn scriptextension_gd_get_method_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetMethodInfo(unsafe{&T(voidptr(inst))})
	method := unsafe{&StringName(args[0])}
	*(&Dictionary(ret)) := v_inst.get_method_info_(method)
}

fn scriptextension_gd_is_tool[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionIsTool(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_tool_()
}

fn scriptextension_gd_is_valid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionIsValid(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_valid_()
}

fn scriptextension_gd_is_abstract[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionIsAbstract(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_abstract_()
}

fn scriptextension_gd_get_language[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetLanguage(unsafe{&T(voidptr(inst))})
	*(&ScriptLanguage(ret)) := v_inst.get_language_()
}

fn scriptextension_gd_has_script_signal[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionHasScriptSignal(unsafe{&T(voidptr(inst))})
	signal := unsafe{&StringName(args[0])}
	*(&bool(ret)) := v_inst.has_script_signal_(signal)
}

fn scriptextension_gd_get_script_signal_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetScriptSignalList(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_script_signal_list_()
}

fn scriptextension_gd_has_property_default_value[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionHasPropertyDefaultValue(unsafe{&T(voidptr(inst))})
	property := unsafe{&StringName(args[0])}
	*(&bool(ret)) := v_inst.has_property_default_value_(property)
}

fn scriptextension_gd_get_property_default_value[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetPropertyDefaultValue(unsafe{&T(voidptr(inst))})
	property := unsafe{&StringName(args[0])}
	*(&Variant(ret)) := v_inst.get_property_default_value_(property)
}

fn scriptextension_gd_update_exports[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionUpdateExports(unsafe{&T(voidptr(inst))})
	v_inst.update_exports_()
}

fn scriptextension_gd_get_script_method_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetScriptMethodList(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_script_method_list_()
}

fn scriptextension_gd_get_script_property_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetScriptPropertyList(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_script_property_list_()
}

fn scriptextension_gd_get_member_line[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetMemberLine(unsafe{&T(voidptr(inst))})
	member := unsafe{&StringName(args[0])}
	*(&i64(ret)) := v_inst.get_member_line_(member)
}

fn scriptextension_gd_get_constants[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetConstants(unsafe{&T(voidptr(inst))})
	*(&Dictionary(ret)) := v_inst.get_constants_()
}

fn scriptextension_gd_get_members[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetMembers(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_members_()
}

fn scriptextension_gd_is_placeholder_fallback_enabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionIsPlaceholderFallbackEnabled(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_placeholder_fallback_enabled_()
}

fn scriptextension_gd_get_rpc_config[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptExtensionGetRpcConfig(unsafe{&T(voidptr(inst))})
	*(&Variant(ret)) := v_inst.get_rpc_config_()
}

fn scriptlanguageextension_gd_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_name_()
}

fn scriptlanguageextension_gd_init[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionInit(unsafe{&T(voidptr(inst))})
	v_inst.init_()
}

fn scriptlanguageextension_gd_get_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetType(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_type_()
}

fn scriptlanguageextension_gd_get_extension[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetExtension(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_extension_()
}

fn scriptlanguageextension_gd_finish[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionFinish(unsafe{&T(voidptr(inst))})
	v_inst.finish_()
}

fn scriptlanguageextension_gd_get_reserved_words[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetReservedWords(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_reserved_words_()
}

fn scriptlanguageextension_gd_is_control_flow_keyword[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionIsControlFlowKeyword(unsafe{&T(voidptr(inst))})
	keyword := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.is_control_flow_keyword_(keyword)
}

fn scriptlanguageextension_gd_get_comment_delimiters[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetCommentDelimiters(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_comment_delimiters_()
}

fn scriptlanguageextension_gd_get_doc_comment_delimiters[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetDocCommentDelimiters(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_doc_comment_delimiters_()
}

fn scriptlanguageextension_gd_get_string_delimiters[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetStringDelimiters(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_string_delimiters_()
}

fn scriptlanguageextension_gd_make_template[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionMakeTemplate(unsafe{&T(voidptr(inst))})
	template := unsafe{&String(args[0])}
	class_name := unsafe{&String(args[1])}
	base_class_name := unsafe{&String(args[2])}
	*(&Script(ret)) := v_inst.make_template_(template, class_name, base_class_name)
}

fn scriptlanguageextension_gd_get_built_in_templates[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetBuiltInTemplates(unsafe{&T(voidptr(inst))})
	object := unsafe{&StringName(args[0])}
	*(&Array(ret)) := v_inst.get_built_in_templates_(object)
}

fn scriptlanguageextension_gd_is_using_templates[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionIsUsingTemplates(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_using_templates_()
}

fn scriptlanguageextension_gd_validate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionValidate(unsafe{&T(voidptr(inst))})
	script := unsafe{&String(args[0])}
	path := unsafe{&String(args[1])}
	validate_functions := unsafe{&bool(args[2])}
	validate_errors := unsafe{&bool(args[3])}
	validate_warnings := unsafe{&bool(args[4])}
	validate_safe_lines := unsafe{&bool(args[5])}
	*(&Dictionary(ret)) := v_inst.validate_(script, path, validate_functions, validate_errors, validate_warnings, validate_safe_lines)
}

fn scriptlanguageextension_gd_validate_path[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionValidatePath(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&String(ret)) := v_inst.validate_path_(path)
}

fn scriptlanguageextension_gd_create_script[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionCreateScript(unsafe{&T(voidptr(inst))})
	*(&Object(ret)) := v_inst.create_script_()
}

fn scriptlanguageextension_gd_has_named_classes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionHasNamedClasses(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_named_classes_()
}

fn scriptlanguageextension_gd_supports_builtin_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionSupportsBuiltinMode(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.supports_builtin_mode_()
}

fn scriptlanguageextension_gd_supports_documentation[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionSupportsDocumentation(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.supports_documentation_()
}

fn scriptlanguageextension_gd_can_inherit_from_file[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionCanInheritFromFile(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_inherit_from_file_()
}

fn scriptlanguageextension_gd_find_function[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionFindFunction(unsafe{&T(voidptr(inst))})
	function := unsafe{&String(args[0])}
	code := unsafe{&String(args[1])}
	*(&i64(ret)) := v_inst.find_function_(function, code)
}

fn scriptlanguageextension_gd_make_function[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionMakeFunction(unsafe{&T(voidptr(inst))})
	class_name := unsafe{&String(args[0])}
	function_name := unsafe{&String(args[1])}
	function_args := unsafe{&PackedStringArray(args[2])}
	*(&String(ret)) := v_inst.make_function_(class_name, function_name, function_args)
}

fn scriptlanguageextension_gd_can_make_function[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionCanMakeFunction(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.can_make_function_()
}

fn scriptlanguageextension_gd_open_in_external_editor[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionOpenInExternalEditor(unsafe{&T(voidptr(inst))})
	script := unsafe{&Script(args[0])}
	line := unsafe{&i64(args[1])}
	column := unsafe{&i64(args[2])}
	*(&GDError(ret)) := v_inst.open_in_external_editor_(script, line, column)
}

fn scriptlanguageextension_gd_overrides_external_editor[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionOverridesExternalEditor(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.overrides_external_editor_()
}

fn scriptlanguageextension_gd_preferred_file_name_casing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionPreferredFileNameCasing(unsafe{&T(voidptr(inst))})
	*(&ScriptLanguageScriptNameCasing(ret)) := v_inst.preferred_file_name_casing_()
}

fn scriptlanguageextension_gd_complete_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionCompleteCode(unsafe{&T(voidptr(inst))})
	code := unsafe{&String(args[0])}
	path := unsafe{&String(args[1])}
	owner := unsafe{&Object(args[2])}
	*(&Dictionary(ret)) := v_inst.complete_code_(code, path, owner)
}

fn scriptlanguageextension_gd_lookup_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionLookupCode(unsafe{&T(voidptr(inst))})
	code := unsafe{&String(args[0])}
	symbol := unsafe{&String(args[1])}
	path := unsafe{&String(args[2])}
	owner := unsafe{&Object(args[3])}
	*(&Dictionary(ret)) := v_inst.lookup_code_(code, symbol, path, owner)
}

fn scriptlanguageextension_gd_auto_indent_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionAutoIndentCode(unsafe{&T(voidptr(inst))})
	code := unsafe{&String(args[0])}
	from_line := unsafe{&i64(args[1])}
	to_line := unsafe{&i64(args[2])}
	*(&String(ret)) := v_inst.auto_indent_code_(code, from_line, to_line)
}

fn scriptlanguageextension_gd_add_global_constant[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionAddGlobalConstant(unsafe{&T(voidptr(inst))})
	name := unsafe{&StringName(args[0])}
	value := unsafe{&Variant(args[1])}
	v_inst.add_global_constant_(name, value)
}

fn scriptlanguageextension_gd_add_named_global_constant[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionAddNamedGlobalConstant(unsafe{&T(voidptr(inst))})
	name := unsafe{&StringName(args[0])}
	value := unsafe{&Variant(args[1])}
	v_inst.add_named_global_constant_(name, value)
}

fn scriptlanguageextension_gd_remove_named_global_constant[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionRemoveNamedGlobalConstant(unsafe{&T(voidptr(inst))})
	name := unsafe{&StringName(args[0])}
	v_inst.remove_named_global_constant_(name)
}

fn scriptlanguageextension_gd_thread_enter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionThreadEnter(unsafe{&T(voidptr(inst))})
	v_inst.thread_enter_()
}

fn scriptlanguageextension_gd_thread_exit[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionThreadExit(unsafe{&T(voidptr(inst))})
	v_inst.thread_exit_()
}

fn scriptlanguageextension_gd_debug_get_error[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetError(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.debug_get_error_()
}

fn scriptlanguageextension_gd_debug_get_stack_level_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetStackLevelCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.debug_get_stack_level_count_()
}

fn scriptlanguageextension_gd_debug_get_stack_level_line[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetStackLevelLine(unsafe{&T(voidptr(inst))})
	level := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.debug_get_stack_level_line_(level)
}

fn scriptlanguageextension_gd_debug_get_stack_level_function[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetStackLevelFunction(unsafe{&T(voidptr(inst))})
	level := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.debug_get_stack_level_function_(level)
}

fn scriptlanguageextension_gd_debug_get_stack_level_source[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetStackLevelSource(unsafe{&T(voidptr(inst))})
	level := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.debug_get_stack_level_source_(level)
}

fn scriptlanguageextension_gd_debug_get_stack_level_locals[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetStackLevelLocals(unsafe{&T(voidptr(inst))})
	level := unsafe{&i64(args[0])}
	max_subitems := unsafe{&i64(args[1])}
	max_depth := unsafe{&i64(args[2])}
	*(&Dictionary(ret)) := v_inst.debug_get_stack_level_locals_(level, max_subitems, max_depth)
}

fn scriptlanguageextension_gd_debug_get_stack_level_members[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetStackLevelMembers(unsafe{&T(voidptr(inst))})
	level := unsafe{&i64(args[0])}
	max_subitems := unsafe{&i64(args[1])}
	max_depth := unsafe{&i64(args[2])}
	*(&Dictionary(ret)) := v_inst.debug_get_stack_level_members_(level, max_subitems, max_depth)
}

fn scriptlanguageextension_gd_debug_get_stack_level_instance[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetStackLevelInstance(unsafe{&T(voidptr(inst))})
	level := unsafe{&i64(args[0])}
	*(&voidptr(ret)) := v_inst.debug_get_stack_level_instance_(level)
}

fn scriptlanguageextension_gd_debug_get_globals[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetGlobals(unsafe{&T(voidptr(inst))})
	max_subitems := unsafe{&i64(args[0])}
	max_depth := unsafe{&i64(args[1])}
	*(&Dictionary(ret)) := v_inst.debug_get_globals_(max_subitems, max_depth)
}

fn scriptlanguageextension_gd_debug_parse_stack_level_expression[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugParseStackLevelExpression(unsafe{&T(voidptr(inst))})
	level := unsafe{&i64(args[0])}
	expression := unsafe{&String(args[1])}
	max_subitems := unsafe{&i64(args[2])}
	max_depth := unsafe{&i64(args[3])}
	*(&String(ret)) := v_inst.debug_parse_stack_level_expression_(level, expression, max_subitems, max_depth)
}

fn scriptlanguageextension_gd_debug_get_current_stack_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionDebugGetCurrentStackInfo(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.debug_get_current_stack_info_()
}

fn scriptlanguageextension_gd_reload_all_scripts[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionReloadAllScripts(unsafe{&T(voidptr(inst))})
	v_inst.reload_all_scripts_()
}

fn scriptlanguageextension_gd_reload_scripts[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionReloadScripts(unsafe{&T(voidptr(inst))})
	scripts := unsafe{&Array(args[0])}
	soft_reload := unsafe{&bool(args[1])}
	v_inst.reload_scripts_(scripts, soft_reload)
}

fn scriptlanguageextension_gd_reload_tool_script[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionReloadToolScript(unsafe{&T(voidptr(inst))})
	script := unsafe{&Script(args[0])}
	soft_reload := unsafe{&bool(args[1])}
	v_inst.reload_tool_script_(script, soft_reload)
}

fn scriptlanguageextension_gd_get_recognized_extensions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetRecognizedExtensions(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_recognized_extensions_()
}

fn scriptlanguageextension_gd_get_public_functions[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetPublicFunctions(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_public_functions_()
}

fn scriptlanguageextension_gd_get_public_constants[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetPublicConstants(unsafe{&T(voidptr(inst))})
	*(&Dictionary(ret)) := v_inst.get_public_constants_()
}

fn scriptlanguageextension_gd_get_public_annotations[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetPublicAnnotations(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_public_annotations_()
}

fn scriptlanguageextension_gd_profiling_start[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionProfilingStart(unsafe{&T(voidptr(inst))})
	v_inst.profiling_start_()
}

fn scriptlanguageextension_gd_profiling_stop[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionProfilingStop(unsafe{&T(voidptr(inst))})
	v_inst.profiling_stop_()
}

fn scriptlanguageextension_gd_profiling_set_save_native_calls[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionProfilingSetSaveNativeCalls(unsafe{&T(voidptr(inst))})
	enable := unsafe{&bool(args[0])}
	v_inst.profiling_set_save_native_calls_(enable)
}

fn scriptlanguageextension_gd_profiling_get_accumulated_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionProfilingGetAccumulatedData(unsafe{&T(voidptr(inst))})
	info_array := unsafe{&&ScriptLanguageExtensionProfilingInfo(args[0])}
	info_max := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.profiling_get_accumulated_data_(info_array, info_max)
}

fn scriptlanguageextension_gd_profiling_get_frame_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionProfilingGetFrameData(unsafe{&T(voidptr(inst))})
	info_array := unsafe{&&ScriptLanguageExtensionProfilingInfo(args[0])}
	info_max := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.profiling_get_frame_data_(info_array, info_max)
}

fn scriptlanguageextension_gd_frame[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionFrame(unsafe{&T(voidptr(inst))})
	v_inst.frame_()
}

fn scriptlanguageextension_gd_handles_global_class_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionHandlesGlobalClassType(unsafe{&T(voidptr(inst))})
	gd_type := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.handles_global_class_type_(gd_type)
}

fn scriptlanguageextension_gd_get_global_class_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IScriptLanguageExtensionGetGlobalClassName(unsafe{&T(voidptr(inst))})
	path := unsafe{&String(args[0])}
	*(&Dictionary(ret)) := v_inst.get_global_class_name_(path)
}

fn skeletonmodification2d_gd_execute[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISkeletonModification2DExecute(unsafe{&T(voidptr(inst))})
	delta := unsafe{&f64(args[0])}
	v_inst.execute_(delta)
}

fn skeletonmodification2d_gd_setup_modification[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISkeletonModification2DSetupModification(unsafe{&T(voidptr(inst))})
	modification_stack := unsafe{&SkeletonModificationStack2D(args[0])}
	v_inst.setup_modification_(modification_stack)
}

fn skeletonmodification2d_gd_draw_editor_gizmo[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISkeletonModification2DDrawEditorGizmo(unsafe{&T(voidptr(inst))})
	v_inst.draw_editor_gizmo_()
}

fn skeletonmodifier3d_gd_process_modification_with_delta[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISkeletonModifier3DProcessModificationWithDelta(unsafe{&T(voidptr(inst))})
	delta := unsafe{&f64(args[0])}
	v_inst.process_modification_with_delta_(delta)
}

fn skeletonmodifier3d_gd_process_modification[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISkeletonModifier3DProcessModification(unsafe{&T(voidptr(inst))})
	v_inst.process_modification_()
}

fn streampeerextension_gd_get_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStreamPeerExtensionGetData(unsafe{&T(voidptr(inst))})
	r_buffer := unsafe{&&u8(args[0])}
	r_bytes := unsafe{&i64(args[1])}
	r_received := unsafe{&&i32(args[2])}
	*(&GDError(ret)) := v_inst.get_data_(r_buffer, r_bytes, r_received)
}

fn streampeerextension_gd_get_partial_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStreamPeerExtensionGetPartialData(unsafe{&T(voidptr(inst))})
	r_buffer := unsafe{&&u8(args[0])}
	r_bytes := unsafe{&i64(args[1])}
	r_received := unsafe{&&i32(args[2])}
	*(&GDError(ret)) := v_inst.get_partial_data_(r_buffer, r_bytes, r_received)
}

fn streampeerextension_gd_put_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStreamPeerExtensionPutData(unsafe{&T(voidptr(inst))})
	p_data := unsafe{&&u8(args[0])}
	p_bytes := unsafe{&i64(args[1])}
	r_sent := unsafe{&&i32(args[2])}
	*(&GDError(ret)) := v_inst.put_data_(p_data, p_bytes, r_sent)
}

fn streampeerextension_gd_put_partial_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStreamPeerExtensionPutPartialData(unsafe{&T(voidptr(inst))})
	p_data := unsafe{&&u8(args[0])}
	p_bytes := unsafe{&i64(args[1])}
	r_sent := unsafe{&&i32(args[2])}
	*(&GDError(ret)) := v_inst.put_partial_data_(p_data, p_bytes, r_sent)
}

fn streampeerextension_gd_get_available_bytes[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStreamPeerExtensionGetAvailableBytes(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_available_bytes_()
}

fn stylebox_gd_draw[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStyleBoxDraw(unsafe{&T(voidptr(inst))})
	to_canvas_item := unsafe{&RID(args[0])}
	rect := unsafe{&Rect2(args[1])}
	v_inst.draw_(to_canvas_item, rect)
}

fn stylebox_gd_get_draw_rect[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStyleBoxGetDrawRect(unsafe{&T(voidptr(inst))})
	rect := unsafe{&Rect2(args[0])}
	*(&Rect2(ret)) := v_inst.get_draw_rect_(rect)
}

fn stylebox_gd_get_minimum_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStyleBoxGetMinimumSize(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_minimum_size_()
}

fn stylebox_gd_test_mask[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IStyleBoxTestMask(unsafe{&T(voidptr(inst))})
	point := unsafe{&Vector2(args[0])}
	rect := unsafe{&Rect2(args[1])}
	*(&bool(ret)) := v_inst.test_mask_(point, rect)
}

fn subviewportcontainer_gd_propagate_input_event[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISubViewportContainerPropagateInputEvent(unsafe{&T(voidptr(inst))})
	event := unsafe{&InputEvent(args[0])}
	*(&bool(ret)) := v_inst.propagate_input_event_(event)
}

fn syntaxhighlighter_gd_get_line_syntax_highlighting[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISyntaxHighlighterGetLineSyntaxHighlighting(unsafe{&T(voidptr(inst))})
	line := unsafe{&i64(args[0])}
	*(&Dictionary(ret)) := v_inst.get_line_syntax_highlighting_(line)
}

fn syntaxhighlighter_gd_clear_highlighting_cache[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISyntaxHighlighterClearHighlightingCache(unsafe{&T(voidptr(inst))})
	v_inst.clear_highlighting_cache_()
}

fn syntaxhighlighter_gd_update_cache[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ISyntaxHighlighterUpdateCache(unsafe{&T(voidptr(inst))})
	v_inst.update_cache_()
}

fn textedit_gd_handle_unicode_input[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextEditHandleUnicodeInput(unsafe{&T(voidptr(inst))})
	unicode_char := unsafe{&i64(args[0])}
	caret_index := unsafe{&i64(args[1])}
	v_inst.handle_unicode_input_(unicode_char, caret_index)
}

fn textedit_gd_backspace[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextEditBackspace(unsafe{&T(voidptr(inst))})
	caret_index := unsafe{&i64(args[0])}
	v_inst.backspace_(caret_index)
}

fn textedit_gd_cut[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextEditCut(unsafe{&T(voidptr(inst))})
	caret_index := unsafe{&i64(args[0])}
	v_inst.cut_(caret_index)
}

fn textedit_gd_copy[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextEditCopy(unsafe{&T(voidptr(inst))})
	caret_index := unsafe{&i64(args[0])}
	v_inst.copy_(caret_index)
}

fn textedit_gd_paste[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextEditPaste(unsafe{&T(voidptr(inst))})
	caret_index := unsafe{&i64(args[0])}
	v_inst.paste_(caret_index)
}

fn textedit_gd_paste_primary_clipboard[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextEditPastePrimaryClipboard(unsafe{&T(voidptr(inst))})
	caret_index := unsafe{&i64(args[0])}
	v_inst.paste_primary_clipboard_(caret_index)
}

fn textserverextension_gd_has_feature[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionHasFeature(unsafe{&T(voidptr(inst))})
	feature := unsafe{&TextServerFeature(args[0])}
	*(&bool(ret)) := v_inst.has_feature_(feature)
}

fn textserverextension_gd_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionGetName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_name_()
}

fn textserverextension_gd_get_features[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionGetFeatures(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_features_()
}

fn textserverextension_gd_free_rid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFreeRid(unsafe{&T(voidptr(inst))})
	rid := unsafe{&RID(args[0])}
	v_inst.free_rid_(rid)
}

fn textserverextension_gd_has[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionHas(unsafe{&T(voidptr(inst))})
	rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.has_(rid)
}

fn textserverextension_gd_load_support_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionLoadSupportData(unsafe{&T(voidptr(inst))})
	filename := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.load_support_data_(filename)
}

fn textserverextension_gd_get_support_data_filename[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionGetSupportDataFilename(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_support_data_filename_()
}

fn textserverextension_gd_get_support_data_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionGetSupportDataInfo(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_support_data_info_()
}

fn textserverextension_gd_save_support_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionSaveSupportData(unsafe{&T(voidptr(inst))})
	filename := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.save_support_data_(filename)
}

fn textserverextension_gd_get_support_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionGetSupportData(unsafe{&T(voidptr(inst))})
	*(&PackedByteArray(ret)) := v_inst.get_support_data_()
}

fn textserverextension_gd_is_locale_right_to_left[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionIsLocaleRightToLeft(unsafe{&T(voidptr(inst))})
	locale := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.is_locale_right_to_left_(locale)
}

fn textserverextension_gd_name_to_tag[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionNameToTag(unsafe{&T(voidptr(inst))})
	name := unsafe{&String(args[0])}
	*(&i64(ret)) := v_inst.name_to_tag_(name)
}

fn textserverextension_gd_tag_to_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionTagToName(unsafe{&T(voidptr(inst))})
	tag := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.tag_to_name_(tag)
}

fn textserverextension_gd_create_font[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionCreateFont(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.create_font_()
}

fn textserverextension_gd_create_font_linked_variation[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionCreateFontLinkedVariation(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&RID(ret)) := v_inst.create_font_linked_variation_(font_rid)
}

fn textserverextension_gd_font_set_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetData(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	data := unsafe{&PackedByteArray(args[1])}
	v_inst.font_set_data_(font_rid, data)
}

fn textserverextension_gd_font_set_data_ptr[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetDataPtr(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	data_ptr := unsafe{&&u8(args[1])}
	data_size := unsafe{&i64(args[2])}
	v_inst.font_set_data_ptr_(font_rid, data_ptr, data_size)
}

fn textserverextension_gd_font_set_face_index[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetFaceIndex(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	face_index := unsafe{&i64(args[1])}
	v_inst.font_set_face_index_(font_rid, face_index)
}

fn textserverextension_gd_font_get_face_index[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetFaceIndex(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.font_get_face_index_(font_rid)
}

fn textserverextension_gd_font_get_face_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetFaceCount(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.font_get_face_count_(font_rid)
}

fn textserverextension_gd_font_set_style[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetStyle(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	style := unsafe{&TextServerFontStyle(args[1])}
	v_inst.font_set_style_(font_rid, style)
}

fn textserverextension_gd_font_get_style[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetStyle(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&TextServerFontStyle(ret)) := v_inst.font_get_style_(font_rid)
}

fn textserverextension_gd_font_set_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetName(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	name := unsafe{&String(args[1])}
	v_inst.font_set_name_(font_rid, name)
}

fn textserverextension_gd_font_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetName(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&String(ret)) := v_inst.font_get_name_(font_rid)
}

fn textserverextension_gd_font_get_ot_name_strings[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetOtNameStrings(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&Dictionary(ret)) := v_inst.font_get_ot_name_strings_(font_rid)
}

fn textserverextension_gd_font_set_style_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetStyleName(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	name_style := unsafe{&String(args[1])}
	v_inst.font_set_style_name_(font_rid, name_style)
}

fn textserverextension_gd_font_get_style_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetStyleName(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&String(ret)) := v_inst.font_get_style_name_(font_rid)
}

fn textserverextension_gd_font_set_weight[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetWeight(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	weight := unsafe{&i64(args[1])}
	v_inst.font_set_weight_(font_rid, weight)
}

fn textserverextension_gd_font_get_weight[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetWeight(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.font_get_weight_(font_rid)
}

fn textserverextension_gd_font_set_stretch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetStretch(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	stretch := unsafe{&i64(args[1])}
	v_inst.font_set_stretch_(font_rid, stretch)
}

fn textserverextension_gd_font_get_stretch[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetStretch(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.font_get_stretch_(font_rid)
}

fn textserverextension_gd_font_set_antialiasing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetAntialiasing(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	antialiasing := unsafe{&TextServerFontAntialiasing(args[1])}
	v_inst.font_set_antialiasing_(font_rid, antialiasing)
}

fn textserverextension_gd_font_get_antialiasing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetAntialiasing(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&TextServerFontAntialiasing(ret)) := v_inst.font_get_antialiasing_(font_rid)
}

fn textserverextension_gd_font_set_disable_embedded_bitmaps[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetDisableEmbeddedBitmaps(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	disable_embedded_bitmaps := unsafe{&bool(args[1])}
	v_inst.font_set_disable_embedded_bitmaps_(font_rid, disable_embedded_bitmaps)
}

fn textserverextension_gd_font_get_disable_embedded_bitmaps[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetDisableEmbeddedBitmaps(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.font_get_disable_embedded_bitmaps_(font_rid)
}

fn textserverextension_gd_font_set_generate_mipmaps[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetGenerateMipmaps(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	generate_mipmaps := unsafe{&bool(args[1])}
	v_inst.font_set_generate_mipmaps_(font_rid, generate_mipmaps)
}

fn textserverextension_gd_font_get_generate_mipmaps[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGenerateMipmaps(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.font_get_generate_mipmaps_(font_rid)
}

fn textserverextension_gd_font_set_multichannel_signed_distance_field[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetMultichannelSignedDistanceField(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	msdf := unsafe{&bool(args[1])}
	v_inst.font_set_multichannel_signed_distance_field_(font_rid, msdf)
}

fn textserverextension_gd_font_is_multichannel_signed_distance_field[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontIsMultichannelSignedDistanceField(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.font_is_multichannel_signed_distance_field_(font_rid)
}

fn textserverextension_gd_font_set_msdf_pixel_range[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetMsdfPixelRange(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	msdf_pixel_range := unsafe{&i64(args[1])}
	v_inst.font_set_msdf_pixel_range_(font_rid, msdf_pixel_range)
}

fn textserverextension_gd_font_get_msdf_pixel_range[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetMsdfPixelRange(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.font_get_msdf_pixel_range_(font_rid)
}

fn textserverextension_gd_font_set_msdf_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetMsdfSize(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	msdf_size := unsafe{&i64(args[1])}
	v_inst.font_set_msdf_size_(font_rid, msdf_size)
}

fn textserverextension_gd_font_get_msdf_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetMsdfSize(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.font_get_msdf_size_(font_rid)
}

fn textserverextension_gd_font_set_fixed_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetFixedSize(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	fixed_size := unsafe{&i64(args[1])}
	v_inst.font_set_fixed_size_(font_rid, fixed_size)
}

fn textserverextension_gd_font_get_fixed_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetFixedSize(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.font_get_fixed_size_(font_rid)
}

fn textserverextension_gd_font_set_fixed_size_scale_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetFixedSizeScaleMode(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	fixed_size_scale_mode := unsafe{&TextServerFixedSizeScaleMode(args[1])}
	v_inst.font_set_fixed_size_scale_mode_(font_rid, fixed_size_scale_mode)
}

fn textserverextension_gd_font_get_fixed_size_scale_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetFixedSizeScaleMode(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&TextServerFixedSizeScaleMode(ret)) := v_inst.font_get_fixed_size_scale_mode_(font_rid)
}

fn textserverextension_gd_font_set_allow_system_fallback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetAllowSystemFallback(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	allow_system_fallback := unsafe{&bool(args[1])}
	v_inst.font_set_allow_system_fallback_(font_rid, allow_system_fallback)
}

fn textserverextension_gd_font_is_allow_system_fallback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontIsAllowSystemFallback(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.font_is_allow_system_fallback_(font_rid)
}

fn textserverextension_gd_font_set_force_autohinter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetForceAutohinter(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	force_autohinter := unsafe{&bool(args[1])}
	v_inst.font_set_force_autohinter_(font_rid, force_autohinter)
}

fn textserverextension_gd_font_is_force_autohinter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontIsForceAutohinter(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.font_is_force_autohinter_(font_rid)
}

fn textserverextension_gd_font_set_modulate_color_glyphs[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetModulateColorGlyphs(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	modulate := unsafe{&bool(args[1])}
	v_inst.font_set_modulate_color_glyphs_(font_rid, modulate)
}

fn textserverextension_gd_font_is_modulate_color_glyphs[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontIsModulateColorGlyphs(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.font_is_modulate_color_glyphs_(font_rid)
}

fn textserverextension_gd_font_set_hinting[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetHinting(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	hinting := unsafe{&TextServerHinting(args[1])}
	v_inst.font_set_hinting_(font_rid, hinting)
}

fn textserverextension_gd_font_get_hinting[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetHinting(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&TextServerHinting(ret)) := v_inst.font_get_hinting_(font_rid)
}

fn textserverextension_gd_font_set_subpixel_positioning[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetSubpixelPositioning(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	subpixel_positioning := unsafe{&TextServerSubpixelPositioning(args[1])}
	v_inst.font_set_subpixel_positioning_(font_rid, subpixel_positioning)
}

fn textserverextension_gd_font_get_subpixel_positioning[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetSubpixelPositioning(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&TextServerSubpixelPositioning(ret)) := v_inst.font_get_subpixel_positioning_(font_rid)
}

fn textserverextension_gd_font_set_keep_rounding_remainders[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetKeepRoundingRemainders(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	keep_rounding_remainders := unsafe{&bool(args[1])}
	v_inst.font_set_keep_rounding_remainders_(font_rid, keep_rounding_remainders)
}

fn textserverextension_gd_font_get_keep_rounding_remainders[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetKeepRoundingRemainders(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.font_get_keep_rounding_remainders_(font_rid)
}

fn textserverextension_gd_font_set_embolden[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetEmbolden(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	strength := unsafe{&f64(args[1])}
	v_inst.font_set_embolden_(font_rid, strength)
}

fn textserverextension_gd_font_get_embolden[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetEmbolden(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.font_get_embolden_(font_rid)
}

fn textserverextension_gd_font_set_spacing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetSpacing(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	spacing := unsafe{&TextServerSpacingType(args[1])}
	value := unsafe{&i64(args[2])}
	v_inst.font_set_spacing_(font_rid, spacing, value)
}

fn textserverextension_gd_font_get_spacing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetSpacing(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	spacing := unsafe{&TextServerSpacingType(args[1])}
	*(&i64(ret)) := v_inst.font_get_spacing_(font_rid, spacing)
}

fn textserverextension_gd_font_set_baseline_offset[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetBaselineOffset(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	baseline_offset := unsafe{&f64(args[1])}
	v_inst.font_set_baseline_offset_(font_rid, baseline_offset)
}

fn textserverextension_gd_font_get_baseline_offset[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetBaselineOffset(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.font_get_baseline_offset_(font_rid)
}

fn textserverextension_gd_font_set_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetTransform(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	transform := unsafe{&Transform2D(args[1])}
	v_inst.font_set_transform_(font_rid, transform)
}

fn textserverextension_gd_font_get_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetTransform(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&Transform2D(ret)) := v_inst.font_get_transform_(font_rid)
}

fn textserverextension_gd_font_set_variation_coordinates[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetVariationCoordinates(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	variation_coordinates := unsafe{&Dictionary(args[1])}
	v_inst.font_set_variation_coordinates_(font_rid, variation_coordinates)
}

fn textserverextension_gd_font_get_variation_coordinates[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetVariationCoordinates(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&Dictionary(ret)) := v_inst.font_get_variation_coordinates_(font_rid)
}

fn textserverextension_gd_font_set_oversampling[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetOversampling(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	oversampling := unsafe{&f64(args[1])}
	v_inst.font_set_oversampling_(font_rid, oversampling)
}

fn textserverextension_gd_font_get_oversampling[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetOversampling(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.font_get_oversampling_(font_rid)
}

fn textserverextension_gd_font_get_size_cache_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetSizeCacheList(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&Array(ret)) := v_inst.font_get_size_cache_list_(font_rid)
}

fn textserverextension_gd_font_clear_size_cache[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontClearSizeCache(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	v_inst.font_clear_size_cache_(font_rid)
}

fn textserverextension_gd_font_remove_size_cache[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRemoveSizeCache(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	v_inst.font_remove_size_cache_(font_rid, size)
}

fn textserverextension_gd_font_set_ascent[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetAscent(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	ascent := unsafe{&f64(args[2])}
	v_inst.font_set_ascent_(font_rid, size, ascent)
}

fn textserverextension_gd_font_get_ascent[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetAscent(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.font_get_ascent_(font_rid, size)
}

fn textserverextension_gd_font_set_descent[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetDescent(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	descent := unsafe{&f64(args[2])}
	v_inst.font_set_descent_(font_rid, size, descent)
}

fn textserverextension_gd_font_get_descent[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetDescent(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.font_get_descent_(font_rid, size)
}

fn textserverextension_gd_font_set_underline_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetUnderlinePosition(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	underline_position := unsafe{&f64(args[2])}
	v_inst.font_set_underline_position_(font_rid, size, underline_position)
}

fn textserverextension_gd_font_get_underline_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetUnderlinePosition(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.font_get_underline_position_(font_rid, size)
}

fn textserverextension_gd_font_set_underline_thickness[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetUnderlineThickness(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	underline_thickness := unsafe{&f64(args[2])}
	v_inst.font_set_underline_thickness_(font_rid, size, underline_thickness)
}

fn textserverextension_gd_font_get_underline_thickness[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetUnderlineThickness(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.font_get_underline_thickness_(font_rid, size)
}

fn textserverextension_gd_font_set_scale[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetScale(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	scale := unsafe{&f64(args[2])}
	v_inst.font_set_scale_(font_rid, size, scale)
}

fn textserverextension_gd_font_get_scale[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetScale(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	*(&f64(ret)) := v_inst.font_get_scale_(font_rid, size)
}

fn textserverextension_gd_font_get_texture_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetTextureCount(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	*(&i64(ret)) := v_inst.font_get_texture_count_(font_rid, size)
}

fn textserverextension_gd_font_clear_textures[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontClearTextures(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	v_inst.font_clear_textures_(font_rid, size)
}

fn textserverextension_gd_font_remove_texture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRemoveTexture(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	texture_index := unsafe{&i64(args[2])}
	v_inst.font_remove_texture_(font_rid, size, texture_index)
}

fn textserverextension_gd_font_set_texture_image[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetTextureImage(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	texture_index := unsafe{&i64(args[2])}
	image := unsafe{&Image(args[3])}
	v_inst.font_set_texture_image_(font_rid, size, texture_index, image)
}

fn textserverextension_gd_font_get_texture_image[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetTextureImage(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	texture_index := unsafe{&i64(args[2])}
	*(&Image(ret)) := v_inst.font_get_texture_image_(font_rid, size, texture_index)
}

fn textserverextension_gd_font_set_texture_offsets[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetTextureOffsets(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	texture_index := unsafe{&i64(args[2])}
	offset := unsafe{&PackedInt32Array(args[3])}
	v_inst.font_set_texture_offsets_(font_rid, size, texture_index, offset)
}

fn textserverextension_gd_font_get_texture_offsets[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetTextureOffsets(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	texture_index := unsafe{&i64(args[2])}
	*(&PackedInt32Array(ret)) := v_inst.font_get_texture_offsets_(font_rid, size, texture_index)
}

fn textserverextension_gd_font_get_glyph_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphList(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	*(&PackedInt32Array(ret)) := v_inst.font_get_glyph_list_(font_rid, size)
}

fn textserverextension_gd_font_clear_glyphs[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontClearGlyphs(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	v_inst.font_clear_glyphs_(font_rid, size)
}

fn textserverextension_gd_font_remove_glyph[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRemoveGlyph(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	v_inst.font_remove_glyph_(font_rid, size, glyph)
}

fn textserverextension_gd_font_get_glyph_advance[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphAdvance(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	glyph := unsafe{&i64(args[2])}
	*(&Vector2(ret)) := v_inst.font_get_glyph_advance_(font_rid, size, glyph)
}

fn textserverextension_gd_font_set_glyph_advance[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetGlyphAdvance(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	glyph := unsafe{&i64(args[2])}
	advance := unsafe{&Vector2(args[3])}
	v_inst.font_set_glyph_advance_(font_rid, size, glyph, advance)
}

fn textserverextension_gd_font_get_glyph_offset[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphOffset(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	*(&Vector2(ret)) := v_inst.font_get_glyph_offset_(font_rid, size, glyph)
}

fn textserverextension_gd_font_set_glyph_offset[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetGlyphOffset(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	offset := unsafe{&Vector2(args[3])}
	v_inst.font_set_glyph_offset_(font_rid, size, glyph, offset)
}

fn textserverextension_gd_font_get_glyph_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphSize(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	*(&Vector2(ret)) := v_inst.font_get_glyph_size_(font_rid, size, glyph)
}

fn textserverextension_gd_font_set_glyph_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetGlyphSize(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	gl_size := unsafe{&Vector2(args[3])}
	v_inst.font_set_glyph_size_(font_rid, size, glyph, gl_size)
}

fn textserverextension_gd_font_get_glyph_uv_rect[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphUvRect(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	*(&Rect2(ret)) := v_inst.font_get_glyph_uv_rect_(font_rid, size, glyph)
}

fn textserverextension_gd_font_set_glyph_uv_rect[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetGlyphUvRect(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	uv_rect := unsafe{&Rect2(args[3])}
	v_inst.font_set_glyph_uv_rect_(font_rid, size, glyph, uv_rect)
}

fn textserverextension_gd_font_get_glyph_texture_idx[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphTextureIdx(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	*(&i64(ret)) := v_inst.font_get_glyph_texture_idx_(font_rid, size, glyph)
}

fn textserverextension_gd_font_set_glyph_texture_idx[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetGlyphTextureIdx(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	texture_idx := unsafe{&i64(args[3])}
	v_inst.font_set_glyph_texture_idx_(font_rid, size, glyph, texture_idx)
}

fn textserverextension_gd_font_get_glyph_texture_rid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphTextureRid(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	*(&RID(ret)) := v_inst.font_get_glyph_texture_rid_(font_rid, size, glyph)
}

fn textserverextension_gd_font_get_glyph_texture_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphTextureSize(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	glyph := unsafe{&i64(args[2])}
	*(&Vector2(ret)) := v_inst.font_get_glyph_texture_size_(font_rid, size, glyph)
}

fn textserverextension_gd_font_get_glyph_contours[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphContours(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	index := unsafe{&i64(args[2])}
	*(&Dictionary(ret)) := v_inst.font_get_glyph_contours_(font_rid, size, index)
}

fn textserverextension_gd_font_get_kerning_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetKerningList(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	*(&Array(ret)) := v_inst.font_get_kerning_list_(font_rid, size)
}

fn textserverextension_gd_font_clear_kerning_map[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontClearKerningMap(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	v_inst.font_clear_kerning_map_(font_rid, size)
}

fn textserverextension_gd_font_remove_kerning[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRemoveKerning(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	glyph_pair := unsafe{&Vector2i(args[2])}
	v_inst.font_remove_kerning_(font_rid, size, glyph_pair)
}

fn textserverextension_gd_font_set_kerning[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetKerning(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	glyph_pair := unsafe{&Vector2i(args[2])}
	kerning := unsafe{&Vector2(args[3])}
	v_inst.font_set_kerning_(font_rid, size, glyph_pair, kerning)
}

fn textserverextension_gd_font_get_kerning[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetKerning(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	glyph_pair := unsafe{&Vector2i(args[2])}
	*(&Vector2(ret)) := v_inst.font_get_kerning_(font_rid, size, glyph_pair)
}

fn textserverextension_gd_font_get_glyph_index[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlyphIndex(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	gd_char := unsafe{&i64(args[2])}
	variation_selector := unsafe{&i64(args[3])}
	*(&i64(ret)) := v_inst.font_get_glyph_index_(font_rid, size, gd_char, variation_selector)
}

fn textserverextension_gd_font_get_char_from_glyph_index[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetCharFromGlyphIndex(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	glyph_index := unsafe{&i64(args[2])}
	*(&i64(ret)) := v_inst.font_get_char_from_glyph_index_(font_rid, size, glyph_index)
}

fn textserverextension_gd_font_has_char[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontHasChar(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	gd_char := unsafe{&i64(args[1])}
	*(&bool(ret)) := v_inst.font_has_char_(font_rid, gd_char)
}

fn textserverextension_gd_font_get_supported_chars[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetSupportedChars(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&String(ret)) := v_inst.font_get_supported_chars_(font_rid)
}

fn textserverextension_gd_font_get_supported_glyphs[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetSupportedGlyphs(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&PackedInt32Array(ret)) := v_inst.font_get_supported_glyphs_(font_rid)
}

fn textserverextension_gd_font_render_range[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRenderRange(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	start := unsafe{&i64(args[2])}
	end := unsafe{&i64(args[3])}
	v_inst.font_render_range_(font_rid, size, start, end)
}

fn textserverextension_gd_font_render_glyph[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRenderGlyph(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	size := unsafe{&Vector2i(args[1])}
	index := unsafe{&i64(args[2])}
	v_inst.font_render_glyph_(font_rid, size, index)
}

fn textserverextension_gd_font_draw_glyph[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontDrawGlyph(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	canvas := unsafe{&RID(args[1])}
	size := unsafe{&i64(args[2])}
	pos := unsafe{&Vector2(args[3])}
	index := unsafe{&i64(args[4])}
	color := unsafe{&Color(args[5])}
	v_inst.font_draw_glyph_(font_rid, canvas, size, pos, index, color)
}

fn textserverextension_gd_font_draw_glyph_outline[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontDrawGlyphOutline(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	canvas := unsafe{&RID(args[1])}
	size := unsafe{&i64(args[2])}
	outline_size := unsafe{&i64(args[3])}
	pos := unsafe{&Vector2(args[4])}
	index := unsafe{&i64(args[5])}
	color := unsafe{&Color(args[6])}
	v_inst.font_draw_glyph_outline_(font_rid, canvas, size, outline_size, pos, index, color)
}

fn textserverextension_gd_font_is_language_supported[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontIsLanguageSupported(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	language := unsafe{&String(args[1])}
	*(&bool(ret)) := v_inst.font_is_language_supported_(font_rid, language)
}

fn textserverextension_gd_font_set_language_support_override[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetLanguageSupportOverride(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	language := unsafe{&String(args[1])}
	supported := unsafe{&bool(args[2])}
	v_inst.font_set_language_support_override_(font_rid, language, supported)
}

fn textserverextension_gd_font_get_language_support_override[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetLanguageSupportOverride(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	language := unsafe{&String(args[1])}
	*(&bool(ret)) := v_inst.font_get_language_support_override_(font_rid, language)
}

fn textserverextension_gd_font_remove_language_support_override[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRemoveLanguageSupportOverride(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	language := unsafe{&String(args[1])}
	v_inst.font_remove_language_support_override_(font_rid, language)
}

fn textserverextension_gd_font_get_language_support_overrides[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetLanguageSupportOverrides(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&PackedStringArray(ret)) := v_inst.font_get_language_support_overrides_(font_rid)
}

fn textserverextension_gd_font_is_script_supported[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontIsScriptSupported(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	script := unsafe{&String(args[1])}
	*(&bool(ret)) := v_inst.font_is_script_supported_(font_rid, script)
}

fn textserverextension_gd_font_set_script_support_override[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetScriptSupportOverride(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	script := unsafe{&String(args[1])}
	supported := unsafe{&bool(args[2])}
	v_inst.font_set_script_support_override_(font_rid, script, supported)
}

fn textserverextension_gd_font_get_script_support_override[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetScriptSupportOverride(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	script := unsafe{&String(args[1])}
	*(&bool(ret)) := v_inst.font_get_script_support_override_(font_rid, script)
}

fn textserverextension_gd_font_remove_script_support_override[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontRemoveScriptSupportOverride(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	script := unsafe{&String(args[1])}
	v_inst.font_remove_script_support_override_(font_rid, script)
}

fn textserverextension_gd_font_get_script_support_overrides[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetScriptSupportOverrides(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&PackedStringArray(ret)) := v_inst.font_get_script_support_overrides_(font_rid)
}

fn textserverextension_gd_font_set_opentype_feature_overrides[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetOpentypeFeatureOverrides(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	overrides := unsafe{&Dictionary(args[1])}
	v_inst.font_set_opentype_feature_overrides_(font_rid, overrides)
}

fn textserverextension_gd_font_get_opentype_feature_overrides[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetOpentypeFeatureOverrides(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&Dictionary(ret)) := v_inst.font_get_opentype_feature_overrides_(font_rid)
}

fn textserverextension_gd_font_supported_feature_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSupportedFeatureList(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&Dictionary(ret)) := v_inst.font_supported_feature_list_(font_rid)
}

fn textserverextension_gd_font_supported_variation_list[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSupportedVariationList(unsafe{&T(voidptr(inst))})
	font_rid := unsafe{&RID(args[0])}
	*(&Dictionary(ret)) := v_inst.font_supported_variation_list_(font_rid)
}

fn textserverextension_gd_font_get_global_oversampling[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontGetGlobalOversampling(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.font_get_global_oversampling_()
}

fn textserverextension_gd_font_set_global_oversampling[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFontSetGlobalOversampling(unsafe{&T(voidptr(inst))})
	oversampling := unsafe{&f64(args[0])}
	v_inst.font_set_global_oversampling_(oversampling)
}

fn textserverextension_gd_get_hex_code_box_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionGetHexCodeBoxSize(unsafe{&T(voidptr(inst))})
	size := unsafe{&i64(args[0])}
	index := unsafe{&i64(args[1])}
	*(&Vector2(ret)) := v_inst.get_hex_code_box_size_(size, index)
}

fn textserverextension_gd_draw_hex_code_box[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionDrawHexCodeBox(unsafe{&T(voidptr(inst))})
	canvas := unsafe{&RID(args[0])}
	size := unsafe{&i64(args[1])}
	pos := unsafe{&Vector2(args[2])}
	index := unsafe{&i64(args[3])}
	color := unsafe{&Color(args[4])}
	v_inst.draw_hex_code_box_(canvas, size, pos, index, color)
}

fn textserverextension_gd_create_shaped_text[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionCreateShapedText(unsafe{&T(voidptr(inst))})
	direction := unsafe{&TextServerDirection(args[0])}
	orientation := unsafe{&TextServerOrientation(args[1])}
	*(&RID(ret)) := v_inst.create_shaped_text_(direction, orientation)
}

fn textserverextension_gd_shaped_text_clear[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextClear(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	v_inst.shaped_text_clear_(shaped)
}

fn textserverextension_gd_shaped_text_set_direction[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetDirection(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	direction := unsafe{&TextServerDirection(args[1])}
	v_inst.shaped_text_set_direction_(shaped, direction)
}

fn textserverextension_gd_shaped_text_get_direction[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetDirection(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&TextServerDirection(ret)) := v_inst.shaped_text_get_direction_(shaped)
}

fn textserverextension_gd_shaped_text_get_inferred_direction[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetInferredDirection(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&TextServerDirection(ret)) := v_inst.shaped_text_get_inferred_direction_(shaped)
}

fn textserverextension_gd_shaped_text_set_bidi_override[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetBidiOverride(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	override := unsafe{&Array(args[1])}
	v_inst.shaped_text_set_bidi_override_(shaped, override)
}

fn textserverextension_gd_shaped_text_set_custom_punctuation[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetCustomPunctuation(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	punct := unsafe{&String(args[1])}
	v_inst.shaped_text_set_custom_punctuation_(shaped, punct)
}

fn textserverextension_gd_shaped_text_get_custom_punctuation[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetCustomPunctuation(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&String(ret)) := v_inst.shaped_text_get_custom_punctuation_(shaped)
}

fn textserverextension_gd_shaped_text_set_custom_ellipsis[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetCustomEllipsis(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	gd_char := unsafe{&i64(args[1])}
	v_inst.shaped_text_set_custom_ellipsis_(shaped, gd_char)
}

fn textserverextension_gd_shaped_text_get_custom_ellipsis[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetCustomEllipsis(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.shaped_text_get_custom_ellipsis_(shaped)
}

fn textserverextension_gd_shaped_text_set_orientation[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetOrientation(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	orientation := unsafe{&TextServerOrientation(args[1])}
	v_inst.shaped_text_set_orientation_(shaped, orientation)
}

fn textserverextension_gd_shaped_text_get_orientation[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetOrientation(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&TextServerOrientation(ret)) := v_inst.shaped_text_get_orientation_(shaped)
}

fn textserverextension_gd_shaped_text_set_preserve_invalid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetPreserveInvalid(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	enabled := unsafe{&bool(args[1])}
	v_inst.shaped_text_set_preserve_invalid_(shaped, enabled)
}

fn textserverextension_gd_shaped_text_get_preserve_invalid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetPreserveInvalid(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.shaped_text_get_preserve_invalid_(shaped)
}

fn textserverextension_gd_shaped_text_set_preserve_control[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetPreserveControl(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	enabled := unsafe{&bool(args[1])}
	v_inst.shaped_text_set_preserve_control_(shaped, enabled)
}

fn textserverextension_gd_shaped_text_get_preserve_control[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetPreserveControl(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.shaped_text_get_preserve_control_(shaped)
}

fn textserverextension_gd_shaped_text_set_spacing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSetSpacing(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	spacing := unsafe{&TextServerSpacingType(args[1])}
	value := unsafe{&i64(args[2])}
	v_inst.shaped_text_set_spacing_(shaped, spacing, value)
}

fn textserverextension_gd_shaped_text_get_spacing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetSpacing(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	spacing := unsafe{&TextServerSpacingType(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_get_spacing_(shaped, spacing)
}

fn textserverextension_gd_shaped_text_add_string[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextAddString(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	text := unsafe{&String(args[1])}
	fonts := unsafe{&Array(args[2])}
	size := unsafe{&i64(args[3])}
	opentype_features := unsafe{&Dictionary(args[4])}
	language := unsafe{&String(args[5])}
	meta := unsafe{&Variant(args[6])}
	*(&bool(ret)) := v_inst.shaped_text_add_string_(shaped, text, fonts, size, opentype_features, language, meta)
}

fn textserverextension_gd_shaped_text_add_object[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextAddObject(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	key := unsafe{&Variant(args[1])}
	size := unsafe{&Vector2(args[2])}
	inline_align := unsafe{&InlineAlignment(args[3])}
	length := unsafe{&i64(args[4])}
	baseline := unsafe{&f64(args[5])}
	*(&bool(ret)) := v_inst.shaped_text_add_object_(shaped, key, size, inline_align, length, baseline)
}

fn textserverextension_gd_shaped_text_resize_object[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextResizeObject(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	key := unsafe{&Variant(args[1])}
	size := unsafe{&Vector2(args[2])}
	inline_align := unsafe{&InlineAlignment(args[3])}
	baseline := unsafe{&f64(args[4])}
	*(&bool(ret)) := v_inst.shaped_text_resize_object_(shaped, key, size, inline_align, baseline)
}

fn textserverextension_gd_shaped_get_text[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetText(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&String(ret)) := v_inst.shaped_get_text_(shaped)
}

fn textserverextension_gd_shaped_get_span_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetSpanCount(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.shaped_get_span_count_(shaped)
}

fn textserverextension_gd_shaped_get_span_meta[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetSpanMeta(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&Variant(ret)) := v_inst.shaped_get_span_meta_(shaped, index)
}

fn textserverextension_gd_shaped_get_span_embedded_object[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetSpanEmbeddedObject(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&Variant(ret)) := v_inst.shaped_get_span_embedded_object_(shaped, index)
}

fn textserverextension_gd_shaped_get_span_text[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetSpanText(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&String(ret)) := v_inst.shaped_get_span_text_(shaped, index)
}

fn textserverextension_gd_shaped_get_span_object[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetSpanObject(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&Variant(ret)) := v_inst.shaped_get_span_object_(shaped, index)
}

fn textserverextension_gd_shaped_set_span_update_font[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedSetSpanUpdateFont(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	fonts := unsafe{&Array(args[2])}
	size := unsafe{&i64(args[3])}
	opentype_features := unsafe{&Dictionary(args[4])}
	v_inst.shaped_set_span_update_font_(shaped, index, fonts, size, opentype_features)
}

fn textserverextension_gd_shaped_get_run_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunCount(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.shaped_get_run_count_(shaped)
}

fn textserverextension_gd_shaped_get_run_text[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunText(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&String(ret)) := v_inst.shaped_get_run_text_(shaped, index)
}

fn textserverextension_gd_shaped_get_run_range[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunRange(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&Vector2i(ret)) := v_inst.shaped_get_run_range_(shaped, index)
}

fn textserverextension_gd_shaped_get_run_font_rid[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunFontRid(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&RID(ret)) := v_inst.shaped_get_run_font_rid_(shaped, index)
}

fn textserverextension_gd_shaped_get_run_font_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunFontSize(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.shaped_get_run_font_size_(shaped, index)
}

fn textserverextension_gd_shaped_get_run_language[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunLanguage(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&String(ret)) := v_inst.shaped_get_run_language_(shaped, index)
}

fn textserverextension_gd_shaped_get_run_direction[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunDirection(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&TextServerDirection(ret)) := v_inst.shaped_get_run_direction_(shaped, index)
}

fn textserverextension_gd_shaped_get_run_object[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedGetRunObject(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	index := unsafe{&i64(args[1])}
	*(&Variant(ret)) := v_inst.shaped_get_run_object_(shaped, index)
}

fn textserverextension_gd_shaped_text_substr[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSubstr(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	start := unsafe{&i64(args[1])}
	length := unsafe{&i64(args[2])}
	*(&RID(ret)) := v_inst.shaped_text_substr_(shaped, start, length)
}

fn textserverextension_gd_shaped_text_get_parent[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetParent(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&RID(ret)) := v_inst.shaped_text_get_parent_(shaped)
}

fn textserverextension_gd_shaped_text_fit_to_width[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextFitToWidth(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	width := unsafe{&f64(args[1])}
	justification_flags := unsafe{&TextServerJustificationFlag(args[2])}
	*(&f64(ret)) := v_inst.shaped_text_fit_to_width_(shaped, width, justification_flags)
}

fn textserverextension_gd_shaped_text_tab_align[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextTabAlign(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	tab_stops := unsafe{&PackedFloat32Array(args[1])}
	*(&f64(ret)) := v_inst.shaped_text_tab_align_(shaped, tab_stops)
}

fn textserverextension_gd_shaped_text_shape[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextShape(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.shaped_text_shape_(shaped)
}

fn textserverextension_gd_shaped_text_update_breaks[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextUpdateBreaks(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.shaped_text_update_breaks_(shaped)
}

fn textserverextension_gd_shaped_text_update_justification_ops[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextUpdateJustificationOps(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.shaped_text_update_justification_ops_(shaped)
}

fn textserverextension_gd_shaped_text_is_ready[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextIsReady(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.shaped_text_is_ready_(shaped)
}

fn textserverextension_gd_shaped_text_get_glyphs[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetGlyphs(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&&Glyph(ret)) := v_inst.shaped_text_get_glyphs_(shaped)
}

fn textserverextension_gd_shaped_text_sort_logical[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextSortLogical(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&&Glyph(ret)) := v_inst.shaped_text_sort_logical_(shaped)
}

fn textserverextension_gd_shaped_text_get_glyph_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetGlyphCount(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.shaped_text_get_glyph_count_(shaped)
}

fn textserverextension_gd_shaped_text_get_range[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetRange(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&Vector2i(ret)) := v_inst.shaped_text_get_range_(shaped)
}

fn textserverextension_gd_shaped_text_get_line_breaks_adv[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetLineBreaksAdv(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	width := unsafe{&PackedFloat32Array(args[1])}
	start := unsafe{&i64(args[2])}
	once := unsafe{&bool(args[3])}
	break_flags := unsafe{&TextServerLineBreakFlag(args[4])}
	*(&PackedInt32Array(ret)) := v_inst.shaped_text_get_line_breaks_adv_(shaped, width, start, once, break_flags)
}

fn textserverextension_gd_shaped_text_get_line_breaks[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetLineBreaks(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	width := unsafe{&f64(args[1])}
	start := unsafe{&i64(args[2])}
	break_flags := unsafe{&TextServerLineBreakFlag(args[3])}
	*(&PackedInt32Array(ret)) := v_inst.shaped_text_get_line_breaks_(shaped, width, start, break_flags)
}

fn textserverextension_gd_shaped_text_get_word_breaks[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetWordBreaks(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	grapheme_flags := unsafe{&TextServerGraphemeFlag(args[1])}
	skip_grapheme_flags := unsafe{&TextServerGraphemeFlag(args[2])}
	*(&PackedInt32Array(ret)) := v_inst.shaped_text_get_word_breaks_(shaped, grapheme_flags, skip_grapheme_flags)
}

fn textserverextension_gd_shaped_text_get_trim_pos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetTrimPos(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.shaped_text_get_trim_pos_(shaped)
}

fn textserverextension_gd_shaped_text_get_ellipsis_pos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetEllipsisPos(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.shaped_text_get_ellipsis_pos_(shaped)
}

fn textserverextension_gd_shaped_text_get_ellipsis_glyph_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetEllipsisGlyphCount(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&i64(ret)) := v_inst.shaped_text_get_ellipsis_glyph_count_(shaped)
}

fn textserverextension_gd_shaped_text_get_ellipsis_glyphs[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetEllipsisGlyphs(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&&Glyph(ret)) := v_inst.shaped_text_get_ellipsis_glyphs_(shaped)
}

fn textserverextension_gd_shaped_text_overrun_trim_to_width[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextOverrunTrimToWidth(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	width := unsafe{&f64(args[1])}
	trim_flags := unsafe{&TextServerTextOverrunFlag(args[2])}
	v_inst.shaped_text_overrun_trim_to_width_(shaped, width, trim_flags)
}

fn textserverextension_gd_shaped_text_get_objects[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetObjects(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&Array(ret)) := v_inst.shaped_text_get_objects_(shaped)
}

fn textserverextension_gd_shaped_text_get_object_rect[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetObjectRect(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	key := unsafe{&Variant(args[1])}
	*(&Rect2(ret)) := v_inst.shaped_text_get_object_rect_(shaped, key)
}

fn textserverextension_gd_shaped_text_get_object_range[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetObjectRange(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	key := unsafe{&Variant(args[1])}
	*(&Vector2i(ret)) := v_inst.shaped_text_get_object_range_(shaped, key)
}

fn textserverextension_gd_shaped_text_get_object_glyph[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetObjectGlyph(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	key := unsafe{&Variant(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_get_object_glyph_(shaped, key)
}

fn textserverextension_gd_shaped_text_get_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetSize(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&Vector2(ret)) := v_inst.shaped_text_get_size_(shaped)
}

fn textserverextension_gd_shaped_text_get_ascent[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetAscent(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shaped_text_get_ascent_(shaped)
}

fn textserverextension_gd_shaped_text_get_descent[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetDescent(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shaped_text_get_descent_(shaped)
}

fn textserverextension_gd_shaped_text_get_width[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetWidth(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shaped_text_get_width_(shaped)
}

fn textserverextension_gd_shaped_text_get_underline_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetUnderlinePosition(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shaped_text_get_underline_position_(shaped)
}

fn textserverextension_gd_shaped_text_get_underline_thickness[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetUnderlineThickness(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&f64(ret)) := v_inst.shaped_text_get_underline_thickness_(shaped)
}

fn textserverextension_gd_shaped_text_get_dominant_direction_in_range[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetDominantDirectionInRange(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	start := unsafe{&i64(args[1])}
	end := unsafe{&i64(args[2])}
	*(&i64(ret)) := v_inst.shaped_text_get_dominant_direction_in_range_(shaped, start, end)
}

fn textserverextension_gd_shaped_text_get_carets[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetCarets(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	position := unsafe{&i64(args[1])}
	caret := unsafe{&&CaretInfo(args[2])}
	v_inst.shaped_text_get_carets_(shaped, position, caret)
}

fn textserverextension_gd_shaped_text_get_selection[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetSelection(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	start := unsafe{&i64(args[1])}
	end := unsafe{&i64(args[2])}
	*(&PackedVector2Array(ret)) := v_inst.shaped_text_get_selection_(shaped, start, end)
}

fn textserverextension_gd_shaped_text_hit_test_grapheme[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextHitTestGrapheme(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	coord := unsafe{&f64(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_hit_test_grapheme_(shaped, coord)
}

fn textserverextension_gd_shaped_text_hit_test_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextHitTestPosition(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	coord := unsafe{&f64(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_hit_test_position_(shaped, coord)
}

fn textserverextension_gd_shaped_text_draw[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextDraw(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	canvas := unsafe{&RID(args[1])}
	pos := unsafe{&Vector2(args[2])}
	clip_l := unsafe{&f64(args[3])}
	clip_r := unsafe{&f64(args[4])}
	color := unsafe{&Color(args[5])}
	v_inst.shaped_text_draw_(shaped, canvas, pos, clip_l, clip_r, color)
}

fn textserverextension_gd_shaped_text_draw_outline[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextDrawOutline(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	canvas := unsafe{&RID(args[1])}
	pos := unsafe{&Vector2(args[2])}
	clip_l := unsafe{&f64(args[3])}
	clip_r := unsafe{&f64(args[4])}
	outline_size := unsafe{&i64(args[5])}
	color := unsafe{&Color(args[6])}
	v_inst.shaped_text_draw_outline_(shaped, canvas, pos, clip_l, clip_r, outline_size, color)
}

fn textserverextension_gd_shaped_text_get_grapheme_bounds[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetGraphemeBounds(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	pos := unsafe{&i64(args[1])}
	*(&Vector2(ret)) := v_inst.shaped_text_get_grapheme_bounds_(shaped, pos)
}

fn textserverextension_gd_shaped_text_next_grapheme_pos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextNextGraphemePos(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	pos := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_next_grapheme_pos_(shaped, pos)
}

fn textserverextension_gd_shaped_text_prev_grapheme_pos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextPrevGraphemePos(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	pos := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_prev_grapheme_pos_(shaped, pos)
}

fn textserverextension_gd_shaped_text_get_character_breaks[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextGetCharacterBreaks(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	*(&PackedInt32Array(ret)) := v_inst.shaped_text_get_character_breaks_(shaped)
}

fn textserverextension_gd_shaped_text_next_character_pos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextNextCharacterPos(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	pos := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_next_character_pos_(shaped, pos)
}

fn textserverextension_gd_shaped_text_prev_character_pos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextPrevCharacterPos(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	pos := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_prev_character_pos_(shaped, pos)
}

fn textserverextension_gd_shaped_text_closest_character_pos[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionShapedTextClosestCharacterPos(unsafe{&T(voidptr(inst))})
	shaped := unsafe{&RID(args[0])}
	pos := unsafe{&i64(args[1])}
	*(&i64(ret)) := v_inst.shaped_text_closest_character_pos_(shaped, pos)
}

fn textserverextension_gd_format_number[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionFormatNumber(unsafe{&T(voidptr(inst))})
	number := unsafe{&String(args[0])}
	language := unsafe{&String(args[1])}
	*(&String(ret)) := v_inst.format_number_(number, language)
}

fn textserverextension_gd_parse_number[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionParseNumber(unsafe{&T(voidptr(inst))})
	number := unsafe{&String(args[0])}
	language := unsafe{&String(args[1])}
	*(&String(ret)) := v_inst.parse_number_(number, language)
}

fn textserverextension_gd_percent_sign[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionPercentSign(unsafe{&T(voidptr(inst))})
	language := unsafe{&String(args[0])}
	*(&String(ret)) := v_inst.percent_sign_(language)
}

fn textserverextension_gd_strip_diacritics[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionStripDiacritics(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	*(&String(ret)) := v_inst.strip_diacritics_(gd_string)
}

fn textserverextension_gd_is_valid_identifier[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionIsValidIdentifier(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.is_valid_identifier_(gd_string)
}

fn textserverextension_gd_is_valid_letter[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionIsValidLetter(unsafe{&T(voidptr(inst))})
	unicode := unsafe{&i64(args[0])}
	*(&bool(ret)) := v_inst.is_valid_letter_(unicode)
}

fn textserverextension_gd_string_get_word_breaks[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionStringGetWordBreaks(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	language := unsafe{&String(args[1])}
	chars_per_line := unsafe{&i64(args[2])}
	*(&PackedInt32Array(ret)) := v_inst.string_get_word_breaks_(gd_string, language, chars_per_line)
}

fn textserverextension_gd_string_get_character_breaks[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionStringGetCharacterBreaks(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	language := unsafe{&String(args[1])}
	*(&PackedInt32Array(ret)) := v_inst.string_get_character_breaks_(gd_string, language)
}

fn textserverextension_gd_is_confusable[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionIsConfusable(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	dict := unsafe{&PackedStringArray(args[1])}
	*(&i64(ret)) := v_inst.is_confusable_(gd_string, dict)
}

fn textserverextension_gd_spoof_check[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionSpoofCheck(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	*(&bool(ret)) := v_inst.spoof_check_(gd_string)
}

fn textserverextension_gd_string_to_upper[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionStringToUpper(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	language := unsafe{&String(args[1])}
	*(&String(ret)) := v_inst.string_to_upper_(gd_string, language)
}

fn textserverextension_gd_string_to_lower[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionStringToLower(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	language := unsafe{&String(args[1])}
	*(&String(ret)) := v_inst.string_to_lower_(gd_string, language)
}

fn textserverextension_gd_string_to_title[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionStringToTitle(unsafe{&T(voidptr(inst))})
	gd_string := unsafe{&String(args[0])}
	language := unsafe{&String(args[1])}
	*(&String(ret)) := v_inst.string_to_title_(gd_string, language)
}

fn textserverextension_gd_parse_structured_text[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionParseStructuredText(unsafe{&T(voidptr(inst))})
	parser_type := unsafe{&TextServerStructuredTextParser(args[0])}
	gd_args := unsafe{&Array(args[1])}
	text := unsafe{&String(args[2])}
	*(&Array(ret)) := v_inst.parse_structured_text_(parser_type, gd_args, text)
}

fn textserverextension_gd_cleanup[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextServerExtensionCleanup(unsafe{&T(voidptr(inst))})
	v_inst.cleanup_()
}

fn texture2d_gd_get_width[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture2DGetWidth(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_width_()
}

fn texture2d_gd_get_height[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture2DGetHeight(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_height_()
}

fn texture2d_gd_is_pixel_opaque[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture2DIsPixelOpaque(unsafe{&T(voidptr(inst))})
	x := unsafe{&i64(args[0])}
	y := unsafe{&i64(args[1])}
	*(&bool(ret)) := v_inst.is_pixel_opaque_(x, y)
}

fn texture2d_gd_has_alpha[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture2DHasAlpha(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_alpha_()
}

fn texture2d_gd_draw[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture2DDraw(unsafe{&T(voidptr(inst))})
	to_canvas_item := unsafe{&RID(args[0])}
	pos := unsafe{&Vector2(args[1])}
	modulate := unsafe{&Color(args[2])}
	transpose := unsafe{&bool(args[3])}
	v_inst.draw_(to_canvas_item, pos, modulate, transpose)
}

fn texture2d_gd_draw_rect[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture2DDrawRect(unsafe{&T(voidptr(inst))})
	to_canvas_item := unsafe{&RID(args[0])}
	rect := unsafe{&Rect2(args[1])}
	tile := unsafe{&bool(args[2])}
	modulate := unsafe{&Color(args[3])}
	transpose := unsafe{&bool(args[4])}
	v_inst.draw_rect_(to_canvas_item, rect, tile, modulate, transpose)
}

fn texture2d_gd_draw_rect_region[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture2DDrawRectRegion(unsafe{&T(voidptr(inst))})
	to_canvas_item := unsafe{&RID(args[0])}
	rect := unsafe{&Rect2(args[1])}
	src_rect := unsafe{&Rect2(args[2])}
	modulate := unsafe{&Color(args[3])}
	transpose := unsafe{&bool(args[4])}
	clip_uv := unsafe{&bool(args[5])}
	v_inst.draw_rect_region_(to_canvas_item, rect, src_rect, modulate, transpose, clip_uv)
}

fn texture3d_gd_get_format[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture3DGetFormat(unsafe{&T(voidptr(inst))})
	*(&ImageFormat(ret)) := v_inst.get_format_()
}

fn texture3d_gd_get_width[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture3DGetWidth(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_width_()
}

fn texture3d_gd_get_height[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture3DGetHeight(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_height_()
}

fn texture3d_gd_get_depth[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture3DGetDepth(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_depth_()
}

fn texture3d_gd_has_mipmaps[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture3DHasMipmaps(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_mipmaps_()
}

fn texture3d_gd_get_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITexture3DGetData(unsafe{&T(voidptr(inst))})
	*(&Array(ret)) := v_inst.get_data_()
}

fn texturelayered_gd_get_format[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextureLayeredGetFormat(unsafe{&T(voidptr(inst))})
	*(&ImageFormat(ret)) := v_inst.get_format_()
}

fn texturelayered_gd_get_layered_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextureLayeredGetLayeredType(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_layered_type_()
}

fn texturelayered_gd_get_width[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextureLayeredGetWidth(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_width_()
}

fn texturelayered_gd_get_height[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextureLayeredGetHeight(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_height_()
}

fn texturelayered_gd_get_layers[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextureLayeredGetLayers(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_layers_()
}

fn texturelayered_gd_has_mipmaps[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextureLayeredHasMipmaps(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.has_mipmaps_()
}

fn texturelayered_gd_get_layer_data[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITextureLayeredGetLayerData(unsafe{&T(voidptr(inst))})
	layer_index := unsafe{&i64(args[0])}
	*(&Image(ret)) := v_inst.get_layer_data_(layer_index)
}

fn tilemap_gd_use_tile_data_runtime_update[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITileMapUseTileDataRuntimeUpdate(unsafe{&T(voidptr(inst))})
	layer := unsafe{&i64(args[0])}
	coords := unsafe{&Vector2i(args[1])}
	*(&bool(ret)) := v_inst.use_tile_data_runtime_update_(layer, coords)
}

fn tilemap_gd_tile_data_runtime_update[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITileMapTileDataRuntimeUpdate(unsafe{&T(voidptr(inst))})
	layer := unsafe{&i64(args[0])}
	coords := unsafe{&Vector2i(args[1])}
	tile_data := unsafe{&TileData(args[2])}
	v_inst.tile_data_runtime_update_(layer, coords, tile_data)
}

fn tilemaplayer_gd_use_tile_data_runtime_update[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITileMapLayerUseTileDataRuntimeUpdate(unsafe{&T(voidptr(inst))})
	coords := unsafe{&Vector2i(args[0])}
	*(&bool(ret)) := v_inst.use_tile_data_runtime_update_(coords)
}

fn tilemaplayer_gd_tile_data_runtime_update[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITileMapLayerTileDataRuntimeUpdate(unsafe{&T(voidptr(inst))})
	coords := unsafe{&Vector2i(args[0])}
	tile_data := unsafe{&TileData(args[1])}
	v_inst.tile_data_runtime_update_(coords, tile_data)
}

fn tilemaplayer_gd_update_cells[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITileMapLayerUpdateCells(unsafe{&T(voidptr(inst))})
	coords := unsafe{&Array(args[0])}
	forced_cleanup := unsafe{&bool(args[1])}
	v_inst.update_cells_(coords, forced_cleanup)
}

fn translation_gd_get_plural_message[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITranslationGetPluralMessage(unsafe{&T(voidptr(inst))})
	src_message := unsafe{&StringName(args[0])}
	src_plural_message := unsafe{&StringName(args[1])}
	n := unsafe{&i64(args[2])}
	context := unsafe{&StringName(args[3])}
	*(&StringName(ret)) := v_inst.get_plural_message_(src_message, src_plural_message, n, context)
}

fn translation_gd_get_message[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &ITranslationGetMessage(unsafe{&T(voidptr(inst))})
	src_message := unsafe{&StringName(args[0])}
	context := unsafe{&StringName(args[1])}
	*(&StringName(ret)) := v_inst.get_message_(src_message, context)
}

fn videostream_gd_instantiate_playback[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamInstantiatePlayback(unsafe{&T(voidptr(inst))})
	*(&VideoStreamPlayback(ret)) := v_inst.instantiate_playback_()
}

fn videostreamplayback_gd_stop[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackStop(unsafe{&T(voidptr(inst))})
	v_inst.stop_()
}

fn videostreamplayback_gd_play[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackPlay(unsafe{&T(voidptr(inst))})
	v_inst.play_()
}

fn videostreamplayback_gd_is_playing[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackIsPlaying(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_playing_()
}

fn videostreamplayback_gd_set_paused[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackSetPaused(unsafe{&T(voidptr(inst))})
	paused := unsafe{&bool(args[0])}
	v_inst.set_paused_(paused)
}

fn videostreamplayback_gd_is_paused[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackIsPaused(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_paused_()
}

fn videostreamplayback_gd_get_length[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackGetLength(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_length_()
}

fn videostreamplayback_gd_get_playback_position[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackGetPlaybackPosition(unsafe{&T(voidptr(inst))})
	*(&f64(ret)) := v_inst.get_playback_position_()
}

fn videostreamplayback_gd_seek[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackSeek(unsafe{&T(voidptr(inst))})
	time := unsafe{&f64(args[0])}
	v_inst.seek_(time)
}

fn videostreamplayback_gd_set_audio_track[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackSetAudioTrack(unsafe{&T(voidptr(inst))})
	idx := unsafe{&i64(args[0])}
	v_inst.set_audio_track_(idx)
}

fn videostreamplayback_gd_get_texture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackGetTexture(unsafe{&T(voidptr(inst))})
	*(&Texture2D(ret)) := v_inst.get_texture_()
}

fn videostreamplayback_gd_update[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackUpdate(unsafe{&T(voidptr(inst))})
	delta := unsafe{&f64(args[0])}
	v_inst.update_(delta)
}

fn videostreamplayback_gd_get_channels[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackGetChannels(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_channels_()
}

fn videostreamplayback_gd_get_mix_rate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVideoStreamPlaybackGetMixRate(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_mix_rate_()
}

fn visualinstance3d_gd_get_aabb[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualInstance3DGetAabb(unsafe{&T(voidptr(inst))})
	*(&AABB(ret)) := v_inst.get_aabb_()
}

fn visualshadernodecustom_gd_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetName(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_name_()
}

fn visualshadernodecustom_gd_get_description[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetDescription(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_description_()
}

fn visualshadernodecustom_gd_get_category[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetCategory(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_category_()
}

fn visualshadernodecustom_gd_get_return_icon_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetReturnIconType(unsafe{&T(voidptr(inst))})
	*(&VisualShaderNodePortType(ret)) := v_inst.get_return_icon_type_()
}

fn visualshadernodecustom_gd_get_input_port_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetInputPortCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_input_port_count_()
}

fn visualshadernodecustom_gd_get_input_port_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetInputPortType(unsafe{&T(voidptr(inst))})
	port := unsafe{&i64(args[0])}
	*(&VisualShaderNodePortType(ret)) := v_inst.get_input_port_type_(port)
}

fn visualshadernodecustom_gd_get_input_port_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetInputPortName(unsafe{&T(voidptr(inst))})
	port := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.get_input_port_name_(port)
}

fn visualshadernodecustom_gd_get_input_port_default_value[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetInputPortDefaultValue(unsafe{&T(voidptr(inst))})
	port := unsafe{&i64(args[0])}
	*(&Variant(ret)) := v_inst.get_input_port_default_value_(port)
}

fn visualshadernodecustom_gd_get_default_input_port[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetDefaultInputPort(unsafe{&T(voidptr(inst))})
	gd_type := unsafe{&VisualShaderNodePortType(args[0])}
	*(&i64(ret)) := v_inst.get_default_input_port_(gd_type)
}

fn visualshadernodecustom_gd_get_output_port_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetOutputPortCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_output_port_count_()
}

fn visualshadernodecustom_gd_get_output_port_type[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetOutputPortType(unsafe{&T(voidptr(inst))})
	port := unsafe{&i64(args[0])}
	*(&VisualShaderNodePortType(ret)) := v_inst.get_output_port_type_(port)
}

fn visualshadernodecustom_gd_get_output_port_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetOutputPortName(unsafe{&T(voidptr(inst))})
	port := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.get_output_port_name_(port)
}

fn visualshadernodecustom_gd_get_property_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetPropertyCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_property_count_()
}

fn visualshadernodecustom_gd_get_property_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetPropertyName(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&String(ret)) := v_inst.get_property_name_(index)
}

fn visualshadernodecustom_gd_get_property_default_index[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetPropertyDefaultIndex(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&i64(ret)) := v_inst.get_property_default_index_(index)
}

fn visualshadernodecustom_gd_get_property_options[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetPropertyOptions(unsafe{&T(voidptr(inst))})
	index := unsafe{&i64(args[0])}
	*(&PackedStringArray(ret)) := v_inst.get_property_options_(index)
}

fn visualshadernodecustom_gd_get_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetCode(unsafe{&T(voidptr(inst))})
	input_vars := unsafe{&Array(args[0])}
	output_vars := unsafe{&Array(args[1])}
	mode := unsafe{&ShaderMode(args[2])}
	gd_type := unsafe{&VisualShaderType(args[3])}
	*(&String(ret)) := v_inst.get_code_(input_vars, output_vars, mode, gd_type)
}

fn visualshadernodecustom_gd_get_func_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetFuncCode(unsafe{&T(voidptr(inst))})
	mode := unsafe{&ShaderMode(args[0])}
	gd_type := unsafe{&VisualShaderType(args[1])}
	*(&String(ret)) := v_inst.get_func_code_(mode, gd_type)
}

fn visualshadernodecustom_gd_get_global_code[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomGetGlobalCode(unsafe{&T(voidptr(inst))})
	mode := unsafe{&ShaderMode(args[0])}
	*(&String(ret)) := v_inst.get_global_code_(mode)
}

fn visualshadernodecustom_gd_is_highend[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomIsHighend(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_highend_()
}

fn visualshadernodecustom_gd_is_available[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IVisualShaderNodeCustomIsAvailable(unsafe{&T(voidptr(inst))})
	mode := unsafe{&ShaderMode(args[0])}
	gd_type := unsafe{&VisualShaderType(args[1])}
	*(&bool(ret)) := v_inst.is_available_(mode, gd_type)
}

fn webrtcdatachannelextension_gd_get_packet[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetPacket(unsafe{&T(voidptr(inst))})
	r_buffer := unsafe{&&&u8 (args[0])}
	r_buffer_size := unsafe{&&i32(args[1])}
	*(&GDError(ret)) := v_inst.get_packet_(r_buffer, r_buffer_size)
}

fn webrtcdatachannelextension_gd_put_packet[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionPutPacket(unsafe{&T(voidptr(inst))})
	p_buffer := unsafe{&&u8(args[0])}
	p_buffer_size := unsafe{&i64(args[1])}
	*(&GDError(ret)) := v_inst.put_packet_(p_buffer, p_buffer_size)
}

fn webrtcdatachannelextension_gd_get_available_packet_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetAvailablePacketCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_available_packet_count_()
}

fn webrtcdatachannelextension_gd_get_max_packet_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetMaxPacketSize(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_max_packet_size_()
}

fn webrtcdatachannelextension_gd_poll[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionPoll(unsafe{&T(voidptr(inst))})
	*(&GDError(ret)) := v_inst.poll_()
}

fn webrtcdatachannelextension_gd_close[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionClose(unsafe{&T(voidptr(inst))})
	v_inst.close_()
}

fn webrtcdatachannelextension_gd_set_write_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionSetWriteMode(unsafe{&T(voidptr(inst))})
	p_write_mode := unsafe{&WebRTCDataChannelWriteMode(args[0])}
	v_inst.set_write_mode_(p_write_mode)
}

fn webrtcdatachannelextension_gd_get_write_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetWriteMode(unsafe{&T(voidptr(inst))})
	*(&WebRTCDataChannelWriteMode(ret)) := v_inst.get_write_mode_()
}

fn webrtcdatachannelextension_gd_was_string_packet[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionWasStringPacket(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.was_string_packet_()
}

fn webrtcdatachannelextension_gd_get_ready_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetReadyState(unsafe{&T(voidptr(inst))})
	*(&WebRTCDataChannelChannelState(ret)) := v_inst.get_ready_state_()
}

fn webrtcdatachannelextension_gd_get_label[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetLabel(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_label_()
}

fn webrtcdatachannelextension_gd_is_ordered[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionIsOrdered(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_ordered_()
}

fn webrtcdatachannelextension_gd_get_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetId(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_id_()
}

fn webrtcdatachannelextension_gd_get_max_packet_life_time[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetMaxPacketLifeTime(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_max_packet_life_time_()
}

fn webrtcdatachannelextension_gd_get_max_retransmits[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetMaxRetransmits(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_max_retransmits_()
}

fn webrtcdatachannelextension_gd_get_protocol[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetProtocol(unsafe{&T(voidptr(inst))})
	*(&String(ret)) := v_inst.get_protocol_()
}

fn webrtcdatachannelextension_gd_is_negotiated[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionIsNegotiated(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_negotiated_()
}

fn webrtcdatachannelextension_gd_get_buffered_amount[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCDataChannelExtensionGetBufferedAmount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_buffered_amount_()
}

fn webrtcpeerconnectionextension_gd_get_connection_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionGetConnectionState(unsafe{&T(voidptr(inst))})
	*(&WebRTCPeerConnectionConnectionState(ret)) := v_inst.get_connection_state_()
}

fn webrtcpeerconnectionextension_gd_get_gathering_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionGetGatheringState(unsafe{&T(voidptr(inst))})
	*(&WebRTCPeerConnectionGatheringState(ret)) := v_inst.get_gathering_state_()
}

fn webrtcpeerconnectionextension_gd_get_signaling_state[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionGetSignalingState(unsafe{&T(voidptr(inst))})
	*(&WebRTCPeerConnectionSignalingState(ret)) := v_inst.get_signaling_state_()
}

fn webrtcpeerconnectionextension_gd_initialize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionInitialize(unsafe{&T(voidptr(inst))})
	p_config := unsafe{&Dictionary(args[0])}
	*(&GDError(ret)) := v_inst.initialize_(p_config)
}

fn webrtcpeerconnectionextension_gd_create_data_channel[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionCreateDataChannel(unsafe{&T(voidptr(inst))})
	p_label := unsafe{&String(args[0])}
	p_config := unsafe{&Dictionary(args[1])}
	*(&WebRTCDataChannel(ret)) := v_inst.create_data_channel_(p_label, p_config)
}

fn webrtcpeerconnectionextension_gd_create_offer[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionCreateOffer(unsafe{&T(voidptr(inst))})
	*(&GDError(ret)) := v_inst.create_offer_()
}

fn webrtcpeerconnectionextension_gd_set_remote_description[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionSetRemoteDescription(unsafe{&T(voidptr(inst))})
	p_type := unsafe{&String(args[0])}
	p_sdp := unsafe{&String(args[1])}
	*(&GDError(ret)) := v_inst.set_remote_description_(p_type, p_sdp)
}

fn webrtcpeerconnectionextension_gd_set_local_description[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionSetLocalDescription(unsafe{&T(voidptr(inst))})
	p_type := unsafe{&String(args[0])}
	p_sdp := unsafe{&String(args[1])}
	*(&GDError(ret)) := v_inst.set_local_description_(p_type, p_sdp)
}

fn webrtcpeerconnectionextension_gd_add_ice_candidate[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionAddIceCandidate(unsafe{&T(voidptr(inst))})
	p_sdp_mid_name := unsafe{&String(args[0])}
	p_sdp_mline_index := unsafe{&i64(args[1])}
	p_sdp_name := unsafe{&String(args[2])}
	*(&GDError(ret)) := v_inst.add_ice_candidate_(p_sdp_mid_name, p_sdp_mline_index, p_sdp_name)
}

fn webrtcpeerconnectionextension_gd_poll[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionPoll(unsafe{&T(voidptr(inst))})
	*(&GDError(ret)) := v_inst.poll_()
}

fn webrtcpeerconnectionextension_gd_close[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWebRTCPeerConnectionExtensionClose(unsafe{&T(voidptr(inst))})
	v_inst.close_()
}

fn window_gd_get_contents_minimum_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IWindowGetContentsMinimumSize(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_contents_minimum_size_()
}

fn xrinterfaceextension_gd_get_name[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetName(unsafe{&T(voidptr(inst))})
	*(&StringName(ret)) := v_inst.get_name_()
}

fn xrinterfaceextension_gd_get_capabilities[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetCapabilities(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_capabilities_()
}

fn xrinterfaceextension_gd_is_initialized[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionIsInitialized(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.is_initialized_()
}

fn xrinterfaceextension_gd_initialize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionInitialize(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.initialize_()
}

fn xrinterfaceextension_gd_uninitialize[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionUninitialize(unsafe{&T(voidptr(inst))})
	v_inst.uninitialize_()
}

fn xrinterfaceextension_gd_get_system_info[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetSystemInfo(unsafe{&T(voidptr(inst))})
	*(&Dictionary(ret)) := v_inst.get_system_info_()
}

fn xrinterfaceextension_gd_supports_play_area_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionSupportsPlayAreaMode(unsafe{&T(voidptr(inst))})
	mode := unsafe{&XRInterfacePlayAreaMode(args[0])}
	*(&bool(ret)) := v_inst.supports_play_area_mode_(mode)
}

fn xrinterfaceextension_gd_get_play_area_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetPlayAreaMode(unsafe{&T(voidptr(inst))})
	*(&XRInterfacePlayAreaMode(ret)) := v_inst.get_play_area_mode_()
}

fn xrinterfaceextension_gd_set_play_area_mode[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionSetPlayAreaMode(unsafe{&T(voidptr(inst))})
	mode := unsafe{&XRInterfacePlayAreaMode(args[0])}
	*(&bool(ret)) := v_inst.set_play_area_mode_(mode)
}

fn xrinterfaceextension_gd_get_play_area[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetPlayArea(unsafe{&T(voidptr(inst))})
	*(&PackedVector3Array(ret)) := v_inst.get_play_area_()
}

fn xrinterfaceextension_gd_get_render_target_size[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetRenderTargetSize(unsafe{&T(voidptr(inst))})
	*(&Vector2(ret)) := v_inst.get_render_target_size_()
}

fn xrinterfaceextension_gd_get_view_count[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetViewCount(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_view_count_()
}

fn xrinterfaceextension_gd_get_camera_transform[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetCameraTransform(unsafe{&T(voidptr(inst))})
	*(&Transform3D(ret)) := v_inst.get_camera_transform_()
}

fn xrinterfaceextension_gd_get_transform_for_view[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetTransformForView(unsafe{&T(voidptr(inst))})
	view := unsafe{&i64(args[0])}
	cam_transform := unsafe{&Transform3D(args[1])}
	*(&Transform3D(ret)) := v_inst.get_transform_for_view_(view, cam_transform)
}

fn xrinterfaceextension_gd_get_projection_for_view[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetProjectionForView(unsafe{&T(voidptr(inst))})
	view := unsafe{&i64(args[0])}
	aspect := unsafe{&f64(args[1])}
	z_near := unsafe{&f64(args[2])}
	z_far := unsafe{&f64(args[3])}
	*(&PackedFloat64Array(ret)) := v_inst.get_projection_for_view_(view, aspect, z_near, z_far)
}

fn xrinterfaceextension_gd_get_vrs_texture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetVrsTexture(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_vrs_texture_()
}

fn xrinterfaceextension_gd_process[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionProcess(unsafe{&T(voidptr(inst))})
	v_inst.process_()
}

fn xrinterfaceextension_gd_pre_render[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionPreRender(unsafe{&T(voidptr(inst))})
	v_inst.pre_render_()
}

fn xrinterfaceextension_gd_pre_draw_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionPreDrawViewport(unsafe{&T(voidptr(inst))})
	render_target := unsafe{&RID(args[0])}
	*(&bool(ret)) := v_inst.pre_draw_viewport_(render_target)
}

fn xrinterfaceextension_gd_post_draw_viewport[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionPostDrawViewport(unsafe{&T(voidptr(inst))})
	render_target := unsafe{&RID(args[0])}
	screen_rect := unsafe{&Rect2(args[1])}
	v_inst.post_draw_viewport_(render_target, screen_rect)
}

fn xrinterfaceextension_gd_end_frame[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionEndFrame(unsafe{&T(voidptr(inst))})
	v_inst.end_frame_()
}

fn xrinterfaceextension_gd_get_suggested_tracker_names[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetSuggestedTrackerNames(unsafe{&T(voidptr(inst))})
	*(&PackedStringArray(ret)) := v_inst.get_suggested_tracker_names_()
}

fn xrinterfaceextension_gd_get_suggested_pose_names[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetSuggestedPoseNames(unsafe{&T(voidptr(inst))})
	tracker_name := unsafe{&StringName(args[0])}
	*(&PackedStringArray(ret)) := v_inst.get_suggested_pose_names_(tracker_name)
}

fn xrinterfaceextension_gd_get_tracking_status[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetTrackingStatus(unsafe{&T(voidptr(inst))})
	*(&XRInterfaceTrackingStatus(ret)) := v_inst.get_tracking_status_()
}

fn xrinterfaceextension_gd_trigger_haptic_pulse[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionTriggerHapticPulse(unsafe{&T(voidptr(inst))})
	action_name := unsafe{&String(args[0])}
	tracker_name := unsafe{&StringName(args[1])}
	frequency := unsafe{&f64(args[2])}
	amplitude := unsafe{&f64(args[3])}
	duration_sec := unsafe{&f64(args[4])}
	delay_sec := unsafe{&f64(args[5])}
	v_inst.trigger_haptic_pulse_(action_name, tracker_name, frequency, amplitude, duration_sec, delay_sec)
}

fn xrinterfaceextension_gd_get_anchor_detection_is_enabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetAnchorDetectionIsEnabled(unsafe{&T(voidptr(inst))})
	*(&bool(ret)) := v_inst.get_anchor_detection_is_enabled_()
}

fn xrinterfaceextension_gd_set_anchor_detection_is_enabled[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionSetAnchorDetectionIsEnabled(unsafe{&T(voidptr(inst))})
	enabled := unsafe{&bool(args[0])}
	v_inst.set_anchor_detection_is_enabled_(enabled)
}

fn xrinterfaceextension_gd_get_camera_feed_id[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetCameraFeedId(unsafe{&T(voidptr(inst))})
	*(&i64(ret)) := v_inst.get_camera_feed_id_()
}

fn xrinterfaceextension_gd_get_color_texture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetColorTexture(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_color_texture_()
}

fn xrinterfaceextension_gd_get_depth_texture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetDepthTexture(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_depth_texture_()
}

fn xrinterfaceextension_gd_get_velocity_texture[T] (inst GDExtensionClassInstancePtr, args &GDExtensionConstTypePtr, ret GDExtensionTypePtr) {
	mut v_inst := &IXRInterfaceExtensionGetVelocityTexture(unsafe{&T(voidptr(inst))})
	*(&RID(ret)) := v_inst.get_velocity_texture_()
}
fn register_virtual_methods[T](mut ci ClassInfo) {
	$if T is IAStar2DEstimateCost {{
		// HACK: force function generation
		if false { unsafe { astar2d_gd_estimate_cost[T](nil, nil, nil) } }

		func := astar2d_gd_estimate_cost[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_estimate_cost")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAStar2DComputeCost {{
		// HACK: force function generation
		if false { unsafe { astar2d_gd_compute_cost[T](nil, nil, nil) } }

		func := astar2d_gd_compute_cost[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_compute_cost")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAStar3DEstimateCost {{
		// HACK: force function generation
		if false { unsafe { astar3d_gd_estimate_cost[T](nil, nil, nil) } }

		func := astar3d_gd_estimate_cost[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_estimate_cost")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAStar3DComputeCost {{
		// HACK: force function generation
		if false { unsafe { astar3d_gd_compute_cost[T](nil, nil, nil) } }

		func := astar3d_gd_compute_cost[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_compute_cost")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAStarGrid2DEstimateCost {{
		// HACK: force function generation
		if false { unsafe { astargrid2d_gd_estimate_cost[T](nil, nil, nil) } }

		func := astargrid2d_gd_estimate_cost[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_estimate_cost")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAStarGrid2DComputeCost {{
		// HACK: force function generation
		if false { unsafe { astargrid2d_gd_compute_cost[T](nil, nil, nil) } }

		func := astargrid2d_gd_compute_cost[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_compute_cost")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationMixerPostProcessKeyValue {{
		// HACK: force function generation
		if false { unsafe { animationmixer_gd_post_process_key_value[T](nil, nil, nil) } }

		func := animationmixer_gd_post_process_key_value[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_post_process_key_value")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeGetChildNodes {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_get_child_nodes[T](nil, nil, nil) } }

		func := animationnode_gd_get_child_nodes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_child_nodes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeGetParameterList {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_get_parameter_list[T](nil, nil, nil) } }

		func := animationnode_gd_get_parameter_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_parameter_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeGetChildByName {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_get_child_by_name[T](nil, nil, nil) } }

		func := animationnode_gd_get_child_by_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_child_by_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeGetParameterDefaultValue {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_get_parameter_default_value[T](nil, nil, nil) } }

		func := animationnode_gd_get_parameter_default_value[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_parameter_default_value")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeIsParameterReadOnly {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_is_parameter_read_only[T](nil, nil, nil) } }

		func := animationnode_gd_is_parameter_read_only[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_parameter_read_only")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeProcess {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_process[T](nil, nil, nil) } }

		func := animationnode_gd_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeGetCaption {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_get_caption[T](nil, nil, nil) } }

		func := animationnode_gd_get_caption[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_caption")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeHasFilter {{
		// HACK: force function generation
		if false { unsafe { animationnode_gd_has_filter[T](nil, nil, nil) } }

		func := animationnode_gd_has_filter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_filter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAnimationNodeExtensionProcessAnimationNode {{
		// HACK: force function generation
		if false { unsafe { animationnodeextension_gd_process_animation_node[T](nil, nil, nil) } }

		func := animationnodeextension_gd_process_animation_node[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process_animation_node")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioEffectInstantiate {{
		// HACK: force function generation
		if false { unsafe { audioeffect_gd_instantiate[T](nil, nil, nil) } }

		func := audioeffect_gd_instantiate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_instantiate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioEffectInstanceProcess {{
		// HACK: force function generation
		if false { unsafe { audioeffectinstance_gd_process[T](nil, nil, nil) } }

		func := audioeffectinstance_gd_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioEffectInstanceProcessSilence {{
		// HACK: force function generation
		if false { unsafe { audioeffectinstance_gd_process_silence[T](nil, nil, nil) } }

		func := audioeffectinstance_gd_process_silence[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process_silence")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamInstantiatePlayback {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_instantiate_playback[T](nil, nil, nil) } }

		func := audiostream_gd_instantiate_playback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_instantiate_playback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamGetStreamName {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_get_stream_name[T](nil, nil, nil) } }

		func := audiostream_gd_get_stream_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_stream_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamGetLength {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_get_length[T](nil, nil, nil) } }

		func := audiostream_gd_get_length[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_length")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamIsMonophonic {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_is_monophonic[T](nil, nil, nil) } }

		func := audiostream_gd_is_monophonic[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_monophonic")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamGetBpm {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_get_bpm[T](nil, nil, nil) } }

		func := audiostream_gd_get_bpm[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_bpm")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamGetBeatCount {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_get_beat_count[T](nil, nil, nil) } }

		func := audiostream_gd_get_beat_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_beat_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamGetParameterList {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_get_parameter_list[T](nil, nil, nil) } }

		func := audiostream_gd_get_parameter_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_parameter_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamHasLoop {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_has_loop[T](nil, nil, nil) } }

		func := audiostream_gd_has_loop[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_loop")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamGetBarBeats {{
		// HACK: force function generation
		if false { unsafe { audiostream_gd_get_bar_beats[T](nil, nil, nil) } }

		func := audiostream_gd_get_bar_beats[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_bar_beats")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackStart {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_start[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_start[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_start")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackStop {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_stop[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_stop[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_stop")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackIsPlaying {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_is_playing[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_is_playing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_playing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackGetLoopCount {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_get_loop_count[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_get_loop_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_loop_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackGetPlaybackPosition {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_get_playback_position[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_get_playback_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_playback_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackSeek {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_seek[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_seek[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_seek")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackMix {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_mix[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_mix[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mix")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackTagUsedStreams {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_tag_used_streams[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_tag_used_streams[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_tag_used_streams")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackSetParameter {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_set_parameter[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_set_parameter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_parameter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackGetParameter {{
		// HACK: force function generation
		if false { unsafe { audiostreamplayback_gd_get_parameter[T](nil, nil, nil) } }

		func := audiostreamplayback_gd_get_parameter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_parameter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackResampledMixResampled {{
		// HACK: force function generation
		if false { unsafe { audiostreamplaybackresampled_gd_mix_resampled[T](nil, nil, nil) } }

		func := audiostreamplaybackresampled_gd_mix_resampled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mix_resampled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IAudioStreamPlaybackResampledGetStreamSamplingRate {{
		// HACK: force function generation
		if false { unsafe { audiostreamplaybackresampled_gd_get_stream_sampling_rate[T](nil, nil, nil) } }

		func := audiostreamplaybackresampled_gd_get_stream_sampling_rate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_stream_sampling_rate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IBaseButtonPressed {{
		// HACK: force function generation
		if false { unsafe { basebutton_gd_pressed[T](nil, nil, nil) } }

		func := basebutton_gd_pressed[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pressed")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IBaseButtonToggled {{
		// HACK: force function generation
		if false { unsafe { basebutton_gd_toggled[T](nil, nil, nil) } }

		func := basebutton_gd_toggled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_toggled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICameraFeedActivateFeed {{
		// HACK: force function generation
		if false { unsafe { camerafeed_gd_activate_feed[T](nil, nil, nil) } }

		func := camerafeed_gd_activate_feed[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_activate_feed")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICameraFeedDeactivateFeed {{
		// HACK: force function generation
		if false { unsafe { camerafeed_gd_deactivate_feed[T](nil, nil, nil) } }

		func := camerafeed_gd_deactivate_feed[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_deactivate_feed")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICanvasItemDraw {{
		// HACK: force function generation
		if false { unsafe { canvasitem_gd_draw[T](nil, nil, nil) } }

		func := canvasitem_gd_draw[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICodeEditConfirmCodeCompletion {{
		// HACK: force function generation
		if false { unsafe { codeedit_gd_confirm_code_completion[T](nil, nil, nil) } }

		func := codeedit_gd_confirm_code_completion[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_confirm_code_completion")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICodeEditRequestCodeCompletion {{
		// HACK: force function generation
		if false { unsafe { codeedit_gd_request_code_completion[T](nil, nil, nil) } }

		func := codeedit_gd_request_code_completion[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_request_code_completion")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICodeEditFilterCodeCompletionCandidates {{
		// HACK: force function generation
		if false { unsafe { codeedit_gd_filter_code_completion_candidates[T](nil, nil, nil) } }

		func := codeedit_gd_filter_code_completion_candidates[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_filter_code_completion_candidates")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject2DInputEvent {{
		// HACK: force function generation
		if false { unsafe { collisionobject2d_gd_input_event[T](nil, nil, nil) } }

		func := collisionobject2d_gd_input_event[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_input_event")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject2DMouseEnter {{
		// HACK: force function generation
		if false { unsafe { collisionobject2d_gd_mouse_enter[T](nil, nil, nil) } }

		func := collisionobject2d_gd_mouse_enter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mouse_enter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject2DMouseExit {{
		// HACK: force function generation
		if false { unsafe { collisionobject2d_gd_mouse_exit[T](nil, nil, nil) } }

		func := collisionobject2d_gd_mouse_exit[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mouse_exit")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject2DMouseShapeEnter {{
		// HACK: force function generation
		if false { unsafe { collisionobject2d_gd_mouse_shape_enter[T](nil, nil, nil) } }

		func := collisionobject2d_gd_mouse_shape_enter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mouse_shape_enter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject2DMouseShapeExit {{
		// HACK: force function generation
		if false { unsafe { collisionobject2d_gd_mouse_shape_exit[T](nil, nil, nil) } }

		func := collisionobject2d_gd_mouse_shape_exit[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mouse_shape_exit")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject3DInputEvent {{
		// HACK: force function generation
		if false { unsafe { collisionobject3d_gd_input_event[T](nil, nil, nil) } }

		func := collisionobject3d_gd_input_event[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_input_event")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject3DMouseEnter {{
		// HACK: force function generation
		if false { unsafe { collisionobject3d_gd_mouse_enter[T](nil, nil, nil) } }

		func := collisionobject3d_gd_mouse_enter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mouse_enter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICollisionObject3DMouseExit {{
		// HACK: force function generation
		if false { unsafe { collisionobject3d_gd_mouse_exit[T](nil, nil, nil) } }

		func := collisionobject3d_gd_mouse_exit[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_mouse_exit")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ICompositorEffectRenderCallback {{
		// HACK: force function generation
		if false { unsafe { compositoreffect_gd_render_callback[T](nil, nil, nil) } }

		func := compositoreffect_gd_render_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_render_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IContainerGetAllowedSizeFlagsHorizontal {{
		// HACK: force function generation
		if false { unsafe { container_gd_get_allowed_size_flags_horizontal[T](nil, nil, nil) } }

		func := container_gd_get_allowed_size_flags_horizontal[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_allowed_size_flags_horizontal")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IContainerGetAllowedSizeFlagsVertical {{
		// HACK: force function generation
		if false { unsafe { container_gd_get_allowed_size_flags_vertical[T](nil, nil, nil) } }

		func := container_gd_get_allowed_size_flags_vertical[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_allowed_size_flags_vertical")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlHasPoint {{
		// HACK: force function generation
		if false { unsafe { control_gd_has_point[T](nil, nil, nil) } }

		func := control_gd_has_point[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_point")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlStructuredTextParser {{
		// HACK: force function generation
		if false { unsafe { control_gd_structured_text_parser[T](nil, nil, nil) } }

		func := control_gd_structured_text_parser[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_structured_text_parser")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlGetMinimumSize {{
		// HACK: force function generation
		if false { unsafe { control_gd_get_minimum_size[T](nil, nil, nil) } }

		func := control_gd_get_minimum_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_minimum_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlGetTooltip {{
		// HACK: force function generation
		if false { unsafe { control_gd_get_tooltip[T](nil, nil, nil) } }

		func := control_gd_get_tooltip[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_tooltip")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlGetDragData {{
		// HACK: force function generation
		if false { unsafe { control_gd_get_drag_data[T](nil, nil, nil) } }

		func := control_gd_get_drag_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_drag_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlCanDropData {{
		// HACK: force function generation
		if false { unsafe { control_gd_can_drop_data[T](nil, nil, nil) } }

		func := control_gd_can_drop_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_drop_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlDropData {{
		// HACK: force function generation
		if false { unsafe { control_gd_drop_data[T](nil, nil, nil) } }

		func := control_gd_drop_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_drop_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlMakeCustomTooltip {{
		// HACK: force function generation
		if false { unsafe { control_gd_make_custom_tooltip[T](nil, nil, nil) } }

		func := control_gd_make_custom_tooltip[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_make_custom_tooltip")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlAccessibilityGetContextualInfo {{
		// HACK: force function generation
		if false { unsafe { control_gd_accessibility_get_contextual_info[T](nil, nil, nil) } }

		func := control_gd_accessibility_get_contextual_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_accessibility_get_contextual_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IControlGuiInput {{
		// HACK: force function generation
		if false { unsafe { control_gd_gui_input[T](nil, nil, nil) } }

		func := control_gd_gui_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_gui_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorContextMenuPluginPopupMenu {{
		// HACK: force function generation
		if false { unsafe { editorcontextmenuplugin_gd_popup_menu[T](nil, nil, nil) } }

		func := editorcontextmenuplugin_gd_popup_menu[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_popup_menu")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorDebuggerPluginSetupSession {{
		// HACK: force function generation
		if false { unsafe { editordebuggerplugin_gd_setup_session[T](nil, nil, nil) } }

		func := editordebuggerplugin_gd_setup_session[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_setup_session")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorDebuggerPluginHasCapture {{
		// HACK: force function generation
		if false { unsafe { editordebuggerplugin_gd_has_capture[T](nil, nil, nil) } }

		func := editordebuggerplugin_gd_has_capture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_capture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorDebuggerPluginCapture {{
		// HACK: force function generation
		if false { unsafe { editordebuggerplugin_gd_capture[T](nil, nil, nil) } }

		func := editordebuggerplugin_gd_capture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_capture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorDebuggerPluginGotoScriptLine {{
		// HACK: force function generation
		if false { unsafe { editordebuggerplugin_gd_goto_script_line[T](nil, nil, nil) } }

		func := editordebuggerplugin_gd_goto_script_line[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_goto_script_line")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorDebuggerPluginBreakpointsClearedInTree {{
		// HACK: force function generation
		if false { unsafe { editordebuggerplugin_gd_breakpoints_cleared_in_tree[T](nil, nil, nil) } }

		func := editordebuggerplugin_gd_breakpoints_cleared_in_tree[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_breakpoints_cleared_in_tree")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorDebuggerPluginBreakpointSetInTree {{
		// HACK: force function generation
		if false { unsafe { editordebuggerplugin_gd_breakpoint_set_in_tree[T](nil, nil, nil) } }

		func := editordebuggerplugin_gd_breakpoint_set_in_tree[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_breakpoint_set_in_tree")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetPresetFeatures {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_preset_features[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_preset_features[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_preset_features")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionIsExecutable {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_is_executable[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_is_executable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_executable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetExportOptions {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_export_options[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_export_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionShouldUpdateExportOptions {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_should_update_export_options[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_should_update_export_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_should_update_export_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetExportOptionVisibility {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_export_option_visibility[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_export_option_visibility[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_option_visibility")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetExportOptionWarning {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_export_option_warning[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_export_option_warning[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_option_warning")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetOsName {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_os_name[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_os_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_os_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetName {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_name[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetLogo {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_logo[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_logo[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_logo")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionPollExport {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_poll_export[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_poll_export[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_poll_export")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetOptionsCount {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_options_count[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_options_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_options_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetOptionsTooltip {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_options_tooltip[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_options_tooltip[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_options_tooltip")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetOptionIcon {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_option_icon[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_option_icon[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_option_icon")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetOptionLabel {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_option_label[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_option_label[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_option_label")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetOptionTooltip {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_option_tooltip[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_option_tooltip[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_option_tooltip")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetDeviceArchitecture {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_device_architecture[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_device_architecture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_device_architecture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionCleanup {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_cleanup[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_cleanup[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cleanup")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionRun {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_run[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_run[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_run")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetRunIcon {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_run_icon[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_run_icon[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_run_icon")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionCanExport {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_can_export[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_can_export[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_export")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionHasValidExportConfiguration {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_has_valid_export_configuration[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_has_valid_export_configuration[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_valid_export_configuration")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionHasValidProjectConfiguration {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_has_valid_project_configuration[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_has_valid_project_configuration[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_valid_project_configuration")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetBinaryExtensions {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_binary_extensions[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_binary_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_binary_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionExportProject {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_export_project[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_export_project[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_project")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionExportPack {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_export_pack[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_export_pack[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_pack")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionExportZip {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_export_zip[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_export_zip[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_zip")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionExportPackPatch {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_export_pack_patch[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_export_pack_patch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_pack_patch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionExportZipPatch {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_export_zip_patch[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_export_zip_patch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_zip_patch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetPlatformFeatures {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_platform_features[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_platform_features[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_platform_features")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPlatformExtensionGetDebugProtocol {{
		// HACK: force function generation
		if false { unsafe { editorexportplatformextension_gd_get_debug_protocol[T](nil, nil, nil) } }

		func := editorexportplatformextension_gd_get_debug_protocol[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_debug_protocol")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginExportFile {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_export_file[T](nil, nil, nil) } }

		func := editorexportplugin_gd_export_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginExportBegin {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_export_begin[T](nil, nil, nil) } }

		func := editorexportplugin_gd_export_begin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_begin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginExportEnd {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_export_end[T](nil, nil, nil) } }

		func := editorexportplugin_gd_export_end[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_end")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginBeginCustomizeResources {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_begin_customize_resources[T](nil, nil, nil) } }

		func := editorexportplugin_gd_begin_customize_resources[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_begin_customize_resources")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginCustomizeResource {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_customize_resource[T](nil, nil, nil) } }

		func := editorexportplugin_gd_customize_resource[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_customize_resource")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginBeginCustomizeScenes {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_begin_customize_scenes[T](nil, nil, nil) } }

		func := editorexportplugin_gd_begin_customize_scenes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_begin_customize_scenes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginCustomizeScene {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_customize_scene[T](nil, nil, nil) } }

		func := editorexportplugin_gd_customize_scene[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_customize_scene")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetCustomizationConfigurationHash {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_customization_configuration_hash[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_customization_configuration_hash[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_customization_configuration_hash")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginEndCustomizeScenes {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_end_customize_scenes[T](nil, nil, nil) } }

		func := editorexportplugin_gd_end_customize_scenes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_end_customize_scenes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginEndCustomizeResources {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_end_customize_resources[T](nil, nil, nil) } }

		func := editorexportplugin_gd_end_customize_resources[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_end_customize_resources")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetExportOptions {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_export_options[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_export_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetExportOptionsOverrides {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_export_options_overrides[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_export_options_overrides[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_options_overrides")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginShouldUpdateExportOptions {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_should_update_export_options[T](nil, nil, nil) } }

		func := editorexportplugin_gd_should_update_export_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_should_update_export_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetExportOptionVisibility {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_export_option_visibility[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_export_option_visibility[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_option_visibility")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetExportOptionWarning {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_export_option_warning[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_export_option_warning[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_option_warning")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetExportFeatures {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_export_features[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_export_features[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_export_features")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetName {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_name[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginSupportsPlatform {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_supports_platform[T](nil, nil, nil) } }

		func := editorexportplugin_gd_supports_platform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_supports_platform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetAndroidDependencies {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_android_dependencies[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_android_dependencies[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_android_dependencies")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetAndroidDependenciesMavenRepos {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_android_dependencies_maven_repos[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_android_dependencies_maven_repos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_android_dependencies_maven_repos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetAndroidLibraries {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_android_libraries[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_android_libraries[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_android_libraries")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetAndroidManifestActivityElementContents {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_android_manifest_activity_element_contents[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_android_manifest_activity_element_contents[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_android_manifest_activity_element_contents")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetAndroidManifestApplicationElementContents {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_android_manifest_application_element_contents[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_android_manifest_application_element_contents[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_android_manifest_application_element_contents")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginGetAndroidManifestElementContents {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_get_android_manifest_element_contents[T](nil, nil, nil) } }

		func := editorexportplugin_gd_get_android_manifest_element_contents[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_android_manifest_element_contents")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorExportPluginUpdateAndroidPrebuiltManifest {{
		// HACK: force function generation
		if false { unsafe { editorexportplugin_gd_update_android_prebuilt_manifest[T](nil, nil, nil) } }

		func := editorexportplugin_gd_update_android_prebuilt_manifest[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_update_android_prebuilt_manifest")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorFileSystemImportFormatSupportQueryIsActive {{
		// HACK: force function generation
		if false { unsafe { editorfilesystemimportformatsupportquery_gd_is_active[T](nil, nil, nil) } }

		func := editorfilesystemimportformatsupportquery_gd_is_active[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_active")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorFileSystemImportFormatSupportQueryGetFileExtensions {{
		// HACK: force function generation
		if false { unsafe { editorfilesystemimportformatsupportquery_gd_get_file_extensions[T](nil, nil, nil) } }

		func := editorfilesystemimportformatsupportquery_gd_get_file_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_file_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorFileSystemImportFormatSupportQueryQuery {{
		// HACK: force function generation
		if false { unsafe { editorfilesystemimportformatsupportquery_gd_query[T](nil, nil, nil) } }

		func := editorfilesystemimportformatsupportquery_gd_query[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_query")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetImporterName {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_importer_name[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_importer_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_importer_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetVisibleName {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_visible_name[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_visible_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_visible_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetPresetCount {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_preset_count[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_preset_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_preset_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetPresetName {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_preset_name[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_preset_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_preset_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetRecognizedExtensions {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_recognized_extensions[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_recognized_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_recognized_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetImportOptions {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_import_options[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_import_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_import_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetSaveExtension {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_save_extension[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_save_extension[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_save_extension")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetResourceType {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_resource_type[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_resource_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_resource_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetPriority {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_priority[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetImportOrder {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_import_order[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_import_order[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_import_order")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetFormatVersion {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_format_version[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_format_version[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_format_version")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginGetOptionVisibility {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_get_option_visibility[T](nil, nil, nil) } }

		func := editorimportplugin_gd_get_option_visibility[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_option_visibility")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginImport {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_import[T](nil, nil, nil) } }

		func := editorimportplugin_gd_import[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorImportPluginCanImportThreaded {{
		// HACK: force function generation
		if false { unsafe { editorimportplugin_gd_can_import_threaded[T](nil, nil, nil) } }

		func := editorimportplugin_gd_can_import_threaded[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_import_threaded")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorInspectorPluginCanHandle {{
		// HACK: force function generation
		if false { unsafe { editorinspectorplugin_gd_can_handle[T](nil, nil, nil) } }

		func := editorinspectorplugin_gd_can_handle[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_handle")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorInspectorPluginParseBegin {{
		// HACK: force function generation
		if false { unsafe { editorinspectorplugin_gd_parse_begin[T](nil, nil, nil) } }

		func := editorinspectorplugin_gd_parse_begin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_begin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorInspectorPluginParseCategory {{
		// HACK: force function generation
		if false { unsafe { editorinspectorplugin_gd_parse_category[T](nil, nil, nil) } }

		func := editorinspectorplugin_gd_parse_category[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_category")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorInspectorPluginParseGroup {{
		// HACK: force function generation
		if false { unsafe { editorinspectorplugin_gd_parse_group[T](nil, nil, nil) } }

		func := editorinspectorplugin_gd_parse_group[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_group")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorInspectorPluginParseProperty {{
		// HACK: force function generation
		if false { unsafe { editorinspectorplugin_gd_parse_property[T](nil, nil, nil) } }

		func := editorinspectorplugin_gd_parse_property[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_property")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorInspectorPluginParseEnd {{
		// HACK: force function generation
		if false { unsafe { editorinspectorplugin_gd_parse_end[T](nil, nil, nil) } }

		func := editorinspectorplugin_gd_parse_end[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_end")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoRedraw {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_redraw[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_redraw[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_redraw")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoGetHandleName {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_get_handle_name[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_get_handle_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_handle_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoIsHandleHighlighted {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_is_handle_highlighted[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_is_handle_highlighted[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_handle_highlighted")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoGetHandleValue {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_get_handle_value[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_get_handle_value[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_handle_value")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoBeginHandleAction {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_begin_handle_action[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_begin_handle_action[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_begin_handle_action")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoSetHandle {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_set_handle[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_set_handle[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_handle")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoCommitHandle {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_commit_handle[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_commit_handle[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_commit_handle")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoSubgizmosIntersectRay {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_subgizmos_intersect_ray[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_subgizmos_intersect_ray[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_subgizmos_intersect_ray")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoSubgizmosIntersectFrustum {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_subgizmos_intersect_frustum[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_subgizmos_intersect_frustum[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_subgizmos_intersect_frustum")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoSetSubgizmoTransform {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_set_subgizmo_transform[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_set_subgizmo_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_subgizmo_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoGetSubgizmoTransform {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_get_subgizmo_transform[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_get_subgizmo_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_subgizmo_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoCommitSubgizmos {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmo_gd_commit_subgizmos[T](nil, nil, nil) } }

		func := editornode3dgizmo_gd_commit_subgizmos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_commit_subgizmos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginHasGizmo {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_has_gizmo[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_has_gizmo[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_gizmo")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginCreateGizmo {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_create_gizmo[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_create_gizmo[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_gizmo")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginGetGizmoName {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_get_gizmo_name[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_get_gizmo_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_gizmo_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginGetPriority {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_get_priority[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_get_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginCanBeHidden {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_can_be_hidden[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_can_be_hidden[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_be_hidden")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginIsSelectableWhenHidden {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_is_selectable_when_hidden[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_is_selectable_when_hidden[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_selectable_when_hidden")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginRedraw {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_redraw[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_redraw[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_redraw")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginGetHandleName {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_get_handle_name[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_get_handle_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_handle_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginIsHandleHighlighted {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_is_handle_highlighted[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_is_handle_highlighted[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_handle_highlighted")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginGetHandleValue {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_get_handle_value[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_get_handle_value[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_handle_value")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginBeginHandleAction {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_begin_handle_action[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_begin_handle_action[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_begin_handle_action")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginSetHandle {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_set_handle[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_set_handle[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_handle")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginCommitHandle {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_commit_handle[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_commit_handle[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_commit_handle")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginSubgizmosIntersectRay {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_subgizmos_intersect_ray[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_subgizmos_intersect_ray[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_subgizmos_intersect_ray")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginSubgizmosIntersectFrustum {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_subgizmos_intersect_frustum[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_subgizmos_intersect_frustum[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_subgizmos_intersect_frustum")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginGetSubgizmoTransform {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_get_subgizmo_transform[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_get_subgizmo_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_subgizmo_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginSetSubgizmoTransform {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_set_subgizmo_transform[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_set_subgizmo_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_subgizmo_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorNode3DGizmoPluginCommitSubgizmos {{
		// HACK: force function generation
		if false { unsafe { editornode3dgizmoplugin_gd_commit_subgizmos[T](nil, nil, nil) } }

		func := editornode3dgizmoplugin_gd_commit_subgizmos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_commit_subgizmos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginForwardCanvasGuiInput {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_forward_canvas_gui_input[T](nil, nil, nil) } }

		func := editorplugin_gd_forward_canvas_gui_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_forward_canvas_gui_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginForwardCanvasDrawOverViewport {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_forward_canvas_draw_over_viewport[T](nil, nil, nil) } }

		func := editorplugin_gd_forward_canvas_draw_over_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_forward_canvas_draw_over_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginForwardCanvasForceDrawOverViewport {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_forward_canvas_force_draw_over_viewport[T](nil, nil, nil) } }

		func := editorplugin_gd_forward_canvas_force_draw_over_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_forward_canvas_force_draw_over_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginForward3dGuiInput {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_forward_3d_gui_input[T](nil, nil, nil) } }

		func := editorplugin_gd_forward_3d_gui_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_forward_3d_gui_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginForward3dDrawOverViewport {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_forward_3d_draw_over_viewport[T](nil, nil, nil) } }

		func := editorplugin_gd_forward_3d_draw_over_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_forward_3d_draw_over_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginForward3dForceDrawOverViewport {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_forward_3d_force_draw_over_viewport[T](nil, nil, nil) } }

		func := editorplugin_gd_forward_3d_force_draw_over_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_forward_3d_force_draw_over_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginGetPluginName {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_get_plugin_name[T](nil, nil, nil) } }

		func := editorplugin_gd_get_plugin_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_plugin_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginGetPluginIcon {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_get_plugin_icon[T](nil, nil, nil) } }

		func := editorplugin_gd_get_plugin_icon[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_plugin_icon")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginHasMainScreen {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_has_main_screen[T](nil, nil, nil) } }

		func := editorplugin_gd_has_main_screen[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_main_screen")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginMakeVisible {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_make_visible[T](nil, nil, nil) } }

		func := editorplugin_gd_make_visible[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_make_visible")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginEdit {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_edit[T](nil, nil, nil) } }

		func := editorplugin_gd_edit[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_edit")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginHandles {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_handles[T](nil, nil, nil) } }

		func := editorplugin_gd_handles[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handles")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginGetState {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_get_state[T](nil, nil, nil) } }

		func := editorplugin_gd_get_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginSetState {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_set_state[T](nil, nil, nil) } }

		func := editorplugin_gd_set_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginClear {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_clear[T](nil, nil, nil) } }

		func := editorplugin_gd_clear[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_clear")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginGetUnsavedStatus {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_get_unsaved_status[T](nil, nil, nil) } }

		func := editorplugin_gd_get_unsaved_status[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_unsaved_status")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginSaveExternalData {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_save_external_data[T](nil, nil, nil) } }

		func := editorplugin_gd_save_external_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_save_external_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginApplyChanges {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_apply_changes[T](nil, nil, nil) } }

		func := editorplugin_gd_apply_changes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_changes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginGetBreakpoints {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_get_breakpoints[T](nil, nil, nil) } }

		func := editorplugin_gd_get_breakpoints[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_breakpoints")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginSetWindowLayout {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_set_window_layout[T](nil, nil, nil) } }

		func := editorplugin_gd_set_window_layout[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_window_layout")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginGetWindowLayout {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_get_window_layout[T](nil, nil, nil) } }

		func := editorplugin_gd_get_window_layout[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_window_layout")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginBuild {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_build[T](nil, nil, nil) } }

		func := editorplugin_gd_build[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_build")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginEnablePlugin {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_enable_plugin[T](nil, nil, nil) } }

		func := editorplugin_gd_enable_plugin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_enable_plugin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPluginDisablePlugin {{
		// HACK: force function generation
		if false { unsafe { editorplugin_gd_disable_plugin[T](nil, nil, nil) } }

		func := editorplugin_gd_disable_plugin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_disable_plugin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPropertyUpdateProperty {{
		// HACK: force function generation
		if false { unsafe { editorproperty_gd_update_property[T](nil, nil, nil) } }

		func := editorproperty_gd_update_property[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_update_property")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorPropertySetReadOnly {{
		// HACK: force function generation
		if false { unsafe { editorproperty_gd_set_read_only[T](nil, nil, nil) } }

		func := editorproperty_gd_set_read_only[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_read_only")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourceConversionPluginConvertsTo {{
		// HACK: force function generation
		if false { unsafe { editorresourceconversionplugin_gd_converts_to[T](nil, nil, nil) } }

		func := editorresourceconversionplugin_gd_converts_to[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_converts_to")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourceConversionPluginHandles {{
		// HACK: force function generation
		if false { unsafe { editorresourceconversionplugin_gd_handles[T](nil, nil, nil) } }

		func := editorresourceconversionplugin_gd_handles[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handles")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourceConversionPluginConvert {{
		// HACK: force function generation
		if false { unsafe { editorresourceconversionplugin_gd_convert[T](nil, nil, nil) } }

		func := editorresourceconversionplugin_gd_convert[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_convert")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourcePickerSetCreateOptions {{
		// HACK: force function generation
		if false { unsafe { editorresourcepicker_gd_set_create_options[T](nil, nil, nil) } }

		func := editorresourcepicker_gd_set_create_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_create_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourcePickerHandleMenuSelected {{
		// HACK: force function generation
		if false { unsafe { editorresourcepicker_gd_handle_menu_selected[T](nil, nil, nil) } }

		func := editorresourcepicker_gd_handle_menu_selected[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handle_menu_selected")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourcePreviewGeneratorHandles {{
		// HACK: force function generation
		if false { unsafe { editorresourcepreviewgenerator_gd_handles[T](nil, nil, nil) } }

		func := editorresourcepreviewgenerator_gd_handles[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handles")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourcePreviewGeneratorGenerate {{
		// HACK: force function generation
		if false { unsafe { editorresourcepreviewgenerator_gd_generate[T](nil, nil, nil) } }

		func := editorresourcepreviewgenerator_gd_generate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourcePreviewGeneratorGenerateFromPath {{
		// HACK: force function generation
		if false { unsafe { editorresourcepreviewgenerator_gd_generate_from_path[T](nil, nil, nil) } }

		func := editorresourcepreviewgenerator_gd_generate_from_path[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generate_from_path")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourcePreviewGeneratorGenerateSmallPreviewAutomatically {{
		// HACK: force function generation
		if false { unsafe { editorresourcepreviewgenerator_gd_generate_small_preview_automatically[T](nil, nil, nil) } }

		func := editorresourcepreviewgenerator_gd_generate_small_preview_automatically[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generate_small_preview_automatically")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourcePreviewGeneratorCanGenerateSmallPreview {{
		// HACK: force function generation
		if false { unsafe { editorresourcepreviewgenerator_gd_can_generate_small_preview[T](nil, nil, nil) } }

		func := editorresourcepreviewgenerator_gd_can_generate_small_preview[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_generate_small_preview")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourceTooltipPluginHandles {{
		// HACK: force function generation
		if false { unsafe { editorresourcetooltipplugin_gd_handles[T](nil, nil, nil) } }

		func := editorresourcetooltipplugin_gd_handles[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handles")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorResourceTooltipPluginMakeTooltipForPath {{
		// HACK: force function generation
		if false { unsafe { editorresourcetooltipplugin_gd_make_tooltip_for_path[T](nil, nil, nil) } }

		func := editorresourcetooltipplugin_gd_make_tooltip_for_path[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_make_tooltip_for_path")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorSceneFormatImporterGetExtensions {{
		// HACK: force function generation
		if false { unsafe { editorsceneformatimporter_gd_get_extensions[T](nil, nil, nil) } }

		func := editorsceneformatimporter_gd_get_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorSceneFormatImporterImportScene {{
		// HACK: force function generation
		if false { unsafe { editorsceneformatimporter_gd_import_scene[T](nil, nil, nil) } }

		func := editorsceneformatimporter_gd_import_scene[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import_scene")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorSceneFormatImporterGetImportOptions {{
		// HACK: force function generation
		if false { unsafe { editorsceneformatimporter_gd_get_import_options[T](nil, nil, nil) } }

		func := editorsceneformatimporter_gd_get_import_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_import_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorSceneFormatImporterGetOptionVisibility {{
		// HACK: force function generation
		if false { unsafe { editorsceneformatimporter_gd_get_option_visibility[T](nil, nil, nil) } }

		func := editorsceneformatimporter_gd_get_option_visibility[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_option_visibility")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPostImport {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimport_gd_post_import[T](nil, nil, nil) } }

		func := editorscenepostimport_gd_post_import[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_post_import")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginGetInternalImportOptions {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_get_internal_import_options[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_get_internal_import_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_internal_import_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginGetInternalOptionVisibility {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_get_internal_option_visibility[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_get_internal_option_visibility[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_internal_option_visibility")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginGetInternalOptionUpdateViewRequired {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_get_internal_option_update_view_required[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_get_internal_option_update_view_required[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_internal_option_update_view_required")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginInternalProcess {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_internal_process[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_internal_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_internal_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginGetImportOptions {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_get_import_options[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_get_import_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_import_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginGetOptionVisibility {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_get_option_visibility[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_get_option_visibility[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_option_visibility")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginPreProcess {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_pre_process[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_pre_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pre_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScenePostImportPluginPostProcess {{
		// HACK: force function generation
		if false { unsafe { editorscenepostimportplugin_gd_post_process[T](nil, nil, nil) } }

		func := editorscenepostimportplugin_gd_post_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_post_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorScriptRun {{
		// HACK: force function generation
		if false { unsafe { editorscript_gd_run[T](nil, nil, nil) } }

		func := editorscript_gd_run[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_run")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorSyntaxHighlighterGetName {{
		// HACK: force function generation
		if false { unsafe { editorsyntaxhighlighter_gd_get_name[T](nil, nil, nil) } }

		func := editorsyntaxhighlighter_gd_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorSyntaxHighlighterGetSupportedLanguages {{
		// HACK: force function generation
		if false { unsafe { editorsyntaxhighlighter_gd_get_supported_languages[T](nil, nil, nil) } }

		func := editorsyntaxhighlighter_gd_get_supported_languages[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_supported_languages")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorTranslationParserPluginParseFile {{
		// HACK: force function generation
		if false { unsafe { editortranslationparserplugin_gd_parse_file[T](nil, nil, nil) } }

		func := editortranslationparserplugin_gd_parse_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorTranslationParserPluginGetRecognizedExtensions {{
		// HACK: force function generation
		if false { unsafe { editortranslationparserplugin_gd_get_recognized_extensions[T](nil, nil, nil) } }

		func := editortranslationparserplugin_gd_get_recognized_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_recognized_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceInitialize {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_initialize[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_initialize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_initialize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceSetCredentials {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_set_credentials[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_set_credentials[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_credentials")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetModifiedFilesData {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_modified_files_data[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_modified_files_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_modified_files_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceStageFile {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_stage_file[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_stage_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_stage_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceUnstageFile {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_unstage_file[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_unstage_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_unstage_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceDiscardFile {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_discard_file[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_discard_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_discard_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceCommit {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_commit[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_commit[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_commit")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetDiff {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_diff[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_diff[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_diff")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceShutDown {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_shut_down[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_shut_down[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shut_down")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetVcsName {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_vcs_name[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_vcs_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_vcs_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetPreviousCommits {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_previous_commits[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_previous_commits[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_previous_commits")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetBranchList {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_branch_list[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_branch_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_branch_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetRemotes {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_remotes[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_remotes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_remotes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceCreateBranch {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_create_branch[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_create_branch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_branch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceRemoveBranch {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_remove_branch[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_remove_branch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_remove_branch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceCreateRemote {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_create_remote[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_create_remote[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_remote")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceRemoveRemote {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_remove_remote[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_remove_remote[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_remove_remote")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetCurrentBranchName {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_current_branch_name[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_current_branch_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_current_branch_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceCheckoutBranch {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_checkout_branch[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_checkout_branch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_checkout_branch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfacePull {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_pull[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_pull[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pull")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfacePush {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_push[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_push[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_push")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceFetch {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_fetch[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_fetch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_fetch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEditorVCSInterfaceGetLineDiff {{
		// HACK: force function generation
		if false { unsafe { editorvcsinterface_gd_get_line_diff[T](nil, nil, nil) } }

		func := editorvcsinterface_gd_get_line_diff[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_line_diff")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEngineProfilerToggle {{
		// HACK: force function generation
		if false { unsafe { engineprofiler_gd_toggle[T](nil, nil, nil) } }

		func := engineprofiler_gd_toggle[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_toggle")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEngineProfilerAddFrame {{
		// HACK: force function generation
		if false { unsafe { engineprofiler_gd_add_frame[T](nil, nil, nil) } }

		func := engineprofiler_gd_add_frame[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_frame")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IEngineProfilerTick {{
		// HACK: force function generation
		if false { unsafe { engineprofiler_gd_tick[T](nil, nil, nil) } }

		func := engineprofiler_gd_tick[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_tick")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionImportPreflight {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_import_preflight[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_import_preflight[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import_preflight")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionGetSupportedExtensions {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_get_supported_extensions[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_get_supported_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_supported_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionParseNodeExtensions {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_parse_node_extensions[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_parse_node_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_node_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionParseImageData {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_parse_image_data[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_parse_image_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_image_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionGetImageFileExtension {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_get_image_file_extension[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_get_image_file_extension[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_image_file_extension")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionParseTextureJson {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_parse_texture_json[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_parse_texture_json[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_texture_json")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionImportObjectModelProperty {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_import_object_model_property[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_import_object_model_property[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import_object_model_property")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionImportPostParse {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_import_post_parse[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_import_post_parse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import_post_parse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionImportPreGenerate {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_import_pre_generate[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_import_pre_generate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import_pre_generate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionGenerateSceneNode {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_generate_scene_node[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_generate_scene_node[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generate_scene_node")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionImportNode {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_import_node[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_import_node[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import_node")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionImportPost {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_import_post[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_import_post[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_import_post")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionExportPreflight {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_export_preflight[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_export_preflight[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_preflight")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionConvertSceneNode {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_convert_scene_node[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_convert_scene_node[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_convert_scene_node")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionExportPostConvert {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_export_post_convert[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_export_post_convert[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_post_convert")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionExportPreserialize {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_export_preserialize[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_export_preserialize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_preserialize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionExportObjectModelProperty {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_export_object_model_property[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_export_object_model_property[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_object_model_property")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionGetSaveableImageFormats {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_get_saveable_image_formats[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_get_saveable_image_formats[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_saveable_image_formats")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionSerializeImageToBytes {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_serialize_image_to_bytes[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_serialize_image_to_bytes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_serialize_image_to_bytes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionSaveImageAtPath {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_save_image_at_path[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_save_image_at_path[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_save_image_at_path")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionSerializeTextureJson {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_serialize_texture_json[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_serialize_texture_json[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_serialize_texture_json")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionExportNode {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_export_node[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_export_node[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_node")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGLTFDocumentExtensionExportPost {{
		// HACK: force function generation
		if false { unsafe { gltfdocumentextension_gd_export_post[T](nil, nil, nil) } }

		func := gltfdocumentextension_gd_export_post[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_export_post")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGraphEditIsInInputHotzone {{
		// HACK: force function generation
		if false { unsafe { graphedit_gd_is_in_input_hotzone[T](nil, nil, nil) } }

		func := graphedit_gd_is_in_input_hotzone[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_in_input_hotzone")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGraphEditIsInOutputHotzone {{
		// HACK: force function generation
		if false { unsafe { graphedit_gd_is_in_output_hotzone[T](nil, nil, nil) } }

		func := graphedit_gd_is_in_output_hotzone[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_in_output_hotzone")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGraphEditGetConnectionLine {{
		// HACK: force function generation
		if false { unsafe { graphedit_gd_get_connection_line[T](nil, nil, nil) } }

		func := graphedit_gd_get_connection_line[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_connection_line")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGraphEditIsNodeHoverValid {{
		// HACK: force function generation
		if false { unsafe { graphedit_gd_is_node_hover_valid[T](nil, nil, nil) } }

		func := graphedit_gd_is_node_hover_valid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_node_hover_valid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IGraphNodeDrawPort {{
		// HACK: force function generation
		if false { unsafe { graphnode_gd_draw_port[T](nil, nil, nil) } }

		func := graphnode_gd_draw_port[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw_port")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IImageFormatLoaderExtensionGetRecognizedExtensions {{
		// HACK: force function generation
		if false { unsafe { imageformatloaderextension_gd_get_recognized_extensions[T](nil, nil, nil) } }

		func := imageformatloaderextension_gd_get_recognized_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_recognized_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IImageFormatLoaderExtensionLoadImage {{
		// HACK: force function generation
		if false { unsafe { imageformatloaderextension_gd_load_image[T](nil, nil, nil) } }

		func := imageformatloaderextension_gd_load_image[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_load_image")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMainLoopInitialize {{
		// HACK: force function generation
		if false { unsafe { mainloop_gd_initialize[T](nil, nil, nil) } }

		func := mainloop_gd_initialize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_initialize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMainLoopPhysicsProcess {{
		// HACK: force function generation
		if false { unsafe { mainloop_gd_physics_process[T](nil, nil, nil) } }

		func := mainloop_gd_physics_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_physics_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMainLoopProcess {{
		// HACK: force function generation
		if false { unsafe { mainloop_gd_process[T](nil, nil, nil) } }

		func := mainloop_gd_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMainLoopFinalize {{
		// HACK: force function generation
		if false { unsafe { mainloop_gd_finalize[T](nil, nil, nil) } }

		func := mainloop_gd_finalize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_finalize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMaterialGetShaderRid {{
		// HACK: force function generation
		if false { unsafe { material_gd_get_shader_rid[T](nil, nil, nil) } }

		func := material_gd_get_shader_rid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_shader_rid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMaterialGetShaderMode {{
		// HACK: force function generation
		if false { unsafe { material_gd_get_shader_mode[T](nil, nil, nil) } }

		func := material_gd_get_shader_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_shader_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMaterialCanDoNextPass {{
		// HACK: force function generation
		if false { unsafe { material_gd_can_do_next_pass[T](nil, nil, nil) } }

		func := material_gd_can_do_next_pass[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_do_next_pass")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMaterialCanUseRenderPriority {{
		// HACK: force function generation
		if false { unsafe { material_gd_can_use_render_priority[T](nil, nil, nil) } }

		func := material_gd_can_use_render_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_use_render_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshGetSurfaceCount {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_get_surface_count[T](nil, nil, nil) } }

		func := mesh_gd_get_surface_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_surface_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetArrayLen {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_array_len[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_array_len[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_array_len")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetArrayIndexLen {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_array_index_len[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_array_index_len[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_array_index_len")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetArrays {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_arrays[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_arrays[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_arrays")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetBlendShapeArrays {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_blend_shape_arrays[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_blend_shape_arrays[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_blend_shape_arrays")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetLods {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_lods[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_lods[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_lods")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetFormat {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_format[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_format[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_format")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetPrimitiveType {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_primitive_type[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_primitive_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_primitive_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceSetMaterial {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_set_material[T](nil, nil, nil) } }

		func := mesh_gd_surface_set_material[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_set_material")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSurfaceGetMaterial {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_surface_get_material[T](nil, nil, nil) } }

		func := mesh_gd_surface_get_material[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_surface_get_material")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshGetBlendShapeCount {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_get_blend_shape_count[T](nil, nil, nil) } }

		func := mesh_gd_get_blend_shape_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_blend_shape_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshGetBlendShapeName {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_get_blend_shape_name[T](nil, nil, nil) } }

		func := mesh_gd_get_blend_shape_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_blend_shape_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshSetBlendShapeName {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_set_blend_shape_name[T](nil, nil, nil) } }

		func := mesh_gd_set_blend_shape_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_blend_shape_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMeshGetAabb {{
		// HACK: force function generation
		if false { unsafe { mesh_gd_get_aabb[T](nil, nil, nil) } }

		func := mesh_gd_get_aabb[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_aabb")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMovieWriterGetAudioMixRate {{
		// HACK: force function generation
		if false { unsafe { moviewriter_gd_get_audio_mix_rate[T](nil, nil, nil) } }

		func := moviewriter_gd_get_audio_mix_rate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_audio_mix_rate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMovieWriterGetAudioSpeakerMode {{
		// HACK: force function generation
		if false { unsafe { moviewriter_gd_get_audio_speaker_mode[T](nil, nil, nil) } }

		func := moviewriter_gd_get_audio_speaker_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_audio_speaker_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMovieWriterHandlesFile {{
		// HACK: force function generation
		if false { unsafe { moviewriter_gd_handles_file[T](nil, nil, nil) } }

		func := moviewriter_gd_handles_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handles_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMovieWriterWriteBegin {{
		// HACK: force function generation
		if false { unsafe { moviewriter_gd_write_begin[T](nil, nil, nil) } }

		func := moviewriter_gd_write_begin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_write_begin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMovieWriterWriteFrame {{
		// HACK: force function generation
		if false { unsafe { moviewriter_gd_write_frame[T](nil, nil, nil) } }

		func := moviewriter_gd_write_frame[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_write_frame")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMovieWriterWriteEnd {{
		// HACK: force function generation
		if false { unsafe { moviewriter_gd_write_end[T](nil, nil, nil) } }

		func := moviewriter_gd_write_end[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_write_end")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionPoll {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_poll[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_poll[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_poll")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionSetMultiplayerPeer {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_set_multiplayer_peer[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_set_multiplayer_peer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_multiplayer_peer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionGetMultiplayerPeer {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_get_multiplayer_peer[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_get_multiplayer_peer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_multiplayer_peer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionGetUniqueId {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_get_unique_id[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_get_unique_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_unique_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionGetPeerIds {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_get_peer_ids[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_get_peer_ids[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_peer_ids")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionRpc {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_rpc[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_rpc[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_rpc")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionGetRemoteSenderId {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_get_remote_sender_id[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_get_remote_sender_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_remote_sender_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionObjectConfigurationAdd {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_object_configuration_add[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_object_configuration_add[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_object_configuration_add")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerAPIExtensionObjectConfigurationRemove {{
		// HACK: force function generation
		if false { unsafe { multiplayerapiextension_gd_object_configuration_remove[T](nil, nil, nil) } }

		func := multiplayerapiextension_gd_object_configuration_remove[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_object_configuration_remove")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetPacket {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_packet[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_packet[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_packet")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionPutPacket {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_put_packet[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_put_packet[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_put_packet")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetAvailablePacketCount {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_available_packet_count[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_available_packet_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_available_packet_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetMaxPacketSize {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_max_packet_size[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_max_packet_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_max_packet_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetPacketScript {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_packet_script[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_packet_script[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_packet_script")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionPutPacketScript {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_put_packet_script[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_put_packet_script[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_put_packet_script")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetPacketChannel {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_packet_channel[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_packet_channel[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_packet_channel")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetPacketMode {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_packet_mode[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_packet_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_packet_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionSetTransferChannel {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_set_transfer_channel[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_set_transfer_channel[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_transfer_channel")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetTransferChannel {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_transfer_channel[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_transfer_channel[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_transfer_channel")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionSetTransferMode {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_set_transfer_mode[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_set_transfer_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_transfer_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetTransferMode {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_transfer_mode[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_transfer_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_transfer_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionSetTargetPeer {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_set_target_peer[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_set_target_peer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_target_peer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetPacketPeer {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_packet_peer[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_packet_peer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_packet_peer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionIsServer {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_is_server[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_is_server[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_server")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionPoll {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_poll[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_poll[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_poll")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionClose {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_close[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_close[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_close")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionDisconnectPeer {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_disconnect_peer[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_disconnect_peer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_disconnect_peer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetUniqueId {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_unique_id[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_unique_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_unique_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionSetRefuseNewConnections {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_set_refuse_new_connections[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_set_refuse_new_connections[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_refuse_new_connections")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionIsRefusingNewConnections {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_is_refusing_new_connections[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_is_refusing_new_connections[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_refusing_new_connections")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionIsServerRelaySupported {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_is_server_relay_supported[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_is_server_relay_supported[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_server_relay_supported")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IMultiplayerPeerExtensionGetConnectionStatus {{
		// HACK: force function generation
		if false { unsafe { multiplayerpeerextension_gd_get_connection_status[T](nil, nil, nil) } }

		func := multiplayerpeerextension_gd_get_connection_status[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_connection_status")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeProcess {{
		// HACK: force function generation
		if false { unsafe { node_gd_process[T](nil, nil, nil) } }

		func := node_gd_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodePhysicsProcess {{
		// HACK: force function generation
		if false { unsafe { node_gd_physics_process[T](nil, nil, nil) } }

		func := node_gd_physics_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_physics_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeEnterTree {{
		// HACK: force function generation
		if false { unsafe { node_gd_enter_tree[T](nil, nil, nil) } }

		func := node_gd_enter_tree[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_enter_tree")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeExitTree {{
		// HACK: force function generation
		if false { unsafe { node_gd_exit_tree[T](nil, nil, nil) } }

		func := node_gd_exit_tree[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_exit_tree")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeReady {{
		// HACK: force function generation
		if false { unsafe { node_gd_ready[T](nil, nil, nil) } }

		func := node_gd_ready[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_ready")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeGetConfigurationWarnings {{
		// HACK: force function generation
		if false { unsafe { node_gd_get_configuration_warnings[T](nil, nil, nil) } }

		func := node_gd_get_configuration_warnings[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_configuration_warnings")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeGetAccessibilityConfigurationWarnings {{
		// HACK: force function generation
		if false { unsafe { node_gd_get_accessibility_configuration_warnings[T](nil, nil, nil) } }

		func := node_gd_get_accessibility_configuration_warnings[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_accessibility_configuration_warnings")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeInput {{
		// HACK: force function generation
		if false { unsafe { node_gd_input[T](nil, nil, nil) } }

		func := node_gd_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeShortcutInput {{
		// HACK: force function generation
		if false { unsafe { node_gd_shortcut_input[T](nil, nil, nil) } }

		func := node_gd_shortcut_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shortcut_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeUnhandledInput {{
		// HACK: force function generation
		if false { unsafe { node_gd_unhandled_input[T](nil, nil, nil) } }

		func := node_gd_unhandled_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_unhandled_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeUnhandledKeyInput {{
		// HACK: force function generation
		if false { unsafe { node_gd_unhandled_key_input[T](nil, nil, nil) } }

		func := node_gd_unhandled_key_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_unhandled_key_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeGetFocusedAccessibilityElement {{
		// HACK: force function generation
		if false { unsafe { node_gd_get_focused_accessibility_element[T](nil, nil, nil) } }

		func := node_gd_get_focused_accessibility_element[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_focused_accessibility_element")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is INodeGetAccessibilityContainerName {{
		// HACK: force function generation
		if false { unsafe { node_gd_get_accessibility_container_name[T](nil, nil, nil) } }

		func := node_gd_get_accessibility_container_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_accessibility_container_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRBindingModifierGetDescription {{
		// HACK: force function generation
		if false { unsafe { openxrbindingmodifier_gd_get_description[T](nil, nil, nil) } }

		func := openxrbindingmodifier_gd_get_description[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_description")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRBindingModifierGetIpModification {{
		// HACK: force function generation
		if false { unsafe { openxrbindingmodifier_gd_get_ip_modification[T](nil, nil, nil) } }

		func := openxrbindingmodifier_gd_get_ip_modification[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_ip_modification")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperGetRequestedExtensions {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_get_requested_extensions[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_get_requested_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_requested_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetSystemPropertiesAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_system_properties_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_system_properties_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_system_properties_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetInstanceCreateInfoAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_instance_create_info_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_instance_create_info_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_instance_create_info_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetSessionCreateAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_session_create_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_session_create_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_session_create_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetSwapchainCreateInfoAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_swapchain_create_info_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_swapchain_create_info_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_swapchain_create_info_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetHandJointLocationsAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_hand_joint_locations_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_hand_joint_locations_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_hand_joint_locations_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetProjectionViewsAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_projection_views_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_projection_views_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_projection_views_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetFrameWaitInfoAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_frame_wait_info_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_frame_wait_info_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_frame_wait_info_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetFrameEndInfoAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_frame_end_info_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_frame_end_info_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_frame_end_info_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetViewLocateInfoAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_view_locate_info_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_view_locate_info_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_view_locate_info_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetReferenceSpaceCreateInfoAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_reference_space_create_info_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_reference_space_create_info_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_reference_space_create_info_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperGetCompositionLayerCount {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_get_composition_layer_count[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_get_composition_layer_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_composition_layer_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperGetCompositionLayer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_get_composition_layer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_get_composition_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_composition_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperGetCompositionLayerOrder {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_get_composition_layer_order[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_get_composition_layer_order[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_composition_layer_order")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperGetSuggestedTrackerNames {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_get_suggested_tracker_names[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_get_suggested_tracker_names[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_suggested_tracker_names")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnRegisterMetadata {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_register_metadata[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_register_metadata[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_register_metadata")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnBeforeInstanceCreated {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_before_instance_created[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_before_instance_created[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_before_instance_created")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnInstanceCreated {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_instance_created[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_instance_created[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_instance_created")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnInstanceDestroyed {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_instance_destroyed[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_instance_destroyed[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_instance_destroyed")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnSessionCreated {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_session_created[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_session_created[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_session_created")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnProcess {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_process[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnPreRender {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_pre_render[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_pre_render[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_pre_render")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnMainSwapchainsCreated {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_main_swapchains_created[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_main_swapchains_created[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_main_swapchains_created")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnPreDrawViewport {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_pre_draw_viewport[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_pre_draw_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_pre_draw_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnPostDrawViewport {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_post_draw_viewport[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_post_draw_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_post_draw_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnSessionDestroyed {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_session_destroyed[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_session_destroyed[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_session_destroyed")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateIdle {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_idle[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_idle[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_idle")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateReady {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_ready[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_ready[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_ready")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateSynchronized {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_synchronized[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_synchronized[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_synchronized")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateVisible {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_visible[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_visible[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_visible")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateFocused {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_focused[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_focused[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_focused")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateStopping {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_stopping[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_stopping[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_stopping")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateLossPending {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_loss_pending[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_loss_pending[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_loss_pending")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnStateExiting {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_state_exiting[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_state_exiting[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_state_exiting")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnEventPolled {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_event_polled[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_event_polled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_event_polled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetViewportCompositionLayerAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_viewport_composition_layer_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_viewport_composition_layer_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_viewport_composition_layer_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperGetViewportCompositionLayerExtensionProperties {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_get_viewport_composition_layer_extension_properties[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_get_viewport_composition_layer_extension_properties[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_viewport_composition_layer_extension_properties")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperGetViewportCompositionLayerExtensionPropertyDefaults {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_get_viewport_composition_layer_extension_property_defaults[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_get_viewport_composition_layer_extension_property_defaults[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_viewport_composition_layer_extension_property_defaults")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperOnViewportCompositionLayerDestroyed {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_on_viewport_composition_layer_destroyed[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_on_viewport_composition_layer_destroyed[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_on_viewport_composition_layer_destroyed")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IOpenXRExtensionWrapperSetAndroidSurfaceSwapchainCreateInfoAndGetNextPointer {{
		// HACK: force function generation
		if false { unsafe { openxrextensionwrapper_gd_set_android_surface_swapchain_create_info_and_get_next_pointer[T](nil, nil, nil) } }

		func := openxrextensionwrapper_gd_set_android_surface_swapchain_create_info_and_get_next_pointer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_android_surface_swapchain_create_info_and_get_next_pointer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPacketPeerExtensionGetPacket {{
		// HACK: force function generation
		if false { unsafe { packetpeerextension_gd_get_packet[T](nil, nil, nil) } }

		func := packetpeerextension_gd_get_packet[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_packet")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPacketPeerExtensionPutPacket {{
		// HACK: force function generation
		if false { unsafe { packetpeerextension_gd_put_packet[T](nil, nil, nil) } }

		func := packetpeerextension_gd_put_packet[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_put_packet")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPacketPeerExtensionGetAvailablePacketCount {{
		// HACK: force function generation
		if false { unsafe { packetpeerextension_gd_get_available_packet_count[T](nil, nil, nil) } }

		func := packetpeerextension_gd_get_available_packet_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_available_packet_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPacketPeerExtensionGetMaxPacketSize {{
		// HACK: force function generation
		if false { unsafe { packetpeerextension_gd_get_max_packet_size[T](nil, nil, nil) } }

		func := packetpeerextension_gd_get_max_packet_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_max_packet_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicalBone3DIntegrateForces {{
		// HACK: force function generation
		if false { unsafe { physicalbone3d_gd_integrate_forces[T](nil, nil, nil) } }

		func := physicalbone3d_gd_integrate_forces[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_integrate_forces")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetTotalGravity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_total_gravity[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_total_gravity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_total_gravity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetTotalLinearDamp {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_total_linear_damp[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_total_linear_damp[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_total_linear_damp")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetTotalAngularDamp {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_total_angular_damp[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_total_angular_damp[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_total_angular_damp")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetCenterOfMass {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_center_of_mass[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_center_of_mass[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_center_of_mass")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetCenterOfMassLocal {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_center_of_mass_local[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_center_of_mass_local[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_center_of_mass_local")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetInverseMass {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_inverse_mass[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_inverse_mass[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_inverse_mass")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetInverseInertia {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_inverse_inertia[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_inverse_inertia[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_inverse_inertia")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionSetLinearVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_set_linear_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_set_linear_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_linear_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetLinearVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_linear_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_linear_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_linear_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionSetAngularVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_set_angular_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_set_angular_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_angular_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetAngularVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_angular_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_angular_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_angular_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionSetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_set_transform[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_set_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_transform[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetVelocityAtLocalPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_velocity_at_local_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_velocity_at_local_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_velocity_at_local_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionApplyCentralImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_apply_central_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_apply_central_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_central_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionApplyImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_apply_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_apply_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionApplyTorqueImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_apply_torque_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_apply_torque_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_torque_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionApplyCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_apply_central_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_apply_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionApplyForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_apply_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_apply_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionApplyTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_apply_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_apply_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionAddConstantCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_add_constant_central_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_add_constant_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_constant_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionAddConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_add_constant_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_add_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionAddConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_add_constant_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_add_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionSetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_set_constant_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_set_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_constant_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionSetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_set_constant_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_set_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_constant_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionSetSleepState {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_set_sleep_state[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_set_sleep_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_sleep_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionIsSleeping {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_is_sleeping[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_is_sleeping[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_sleeping")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactCount {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_count[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactLocalPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_local_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_local_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactLocalNormal {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_local_normal[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_local_normal[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_normal")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactLocalShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_local_shape[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_local_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactLocalVelocityAtPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_local_velocity_at_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_local_velocity_at_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_velocity_at_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactCollider {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_collider[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_collider[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactColliderPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_collider_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_collider_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactColliderId {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_collider_id[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_collider_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactColliderObject {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_collider_object[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_collider_object[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_object")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactColliderShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_collider_shape[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_collider_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactColliderVelocityAtPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_collider_velocity_at_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_collider_velocity_at_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_velocity_at_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetContactImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_contact_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_contact_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetStep {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_step[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_step[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_step")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionIntegrateForces {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_integrate_forces[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_integrate_forces[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_integrate_forces")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState2DExtensionGetSpaceState {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate2dextension_gd_get_space_state[T](nil, nil, nil) } }

		func := physicsdirectbodystate2dextension_gd_get_space_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_space_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetTotalGravity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_total_gravity[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_total_gravity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_total_gravity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetTotalLinearDamp {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_total_linear_damp[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_total_linear_damp[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_total_linear_damp")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetTotalAngularDamp {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_total_angular_damp[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_total_angular_damp[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_total_angular_damp")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetCenterOfMass {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_center_of_mass[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_center_of_mass[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_center_of_mass")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetCenterOfMassLocal {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_center_of_mass_local[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_center_of_mass_local[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_center_of_mass_local")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetPrincipalInertiaAxes {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_principal_inertia_axes[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_principal_inertia_axes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_principal_inertia_axes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetInverseMass {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_inverse_mass[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_inverse_mass[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_inverse_mass")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetInverseInertia {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_inverse_inertia[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_inverse_inertia[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_inverse_inertia")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetInverseInertiaTensor {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_inverse_inertia_tensor[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_inverse_inertia_tensor[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_inverse_inertia_tensor")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionSetLinearVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_set_linear_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_set_linear_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_linear_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetLinearVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_linear_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_linear_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_linear_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionSetAngularVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_set_angular_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_set_angular_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_angular_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetAngularVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_angular_velocity[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_angular_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_angular_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionSetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_set_transform[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_set_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_transform[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetVelocityAtLocalPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_velocity_at_local_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_velocity_at_local_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_velocity_at_local_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionApplyCentralImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_apply_central_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_apply_central_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_central_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionApplyImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_apply_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_apply_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionApplyTorqueImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_apply_torque_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_apply_torque_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_torque_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionApplyCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_apply_central_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_apply_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionApplyForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_apply_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_apply_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionApplyTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_apply_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_apply_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_apply_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionAddConstantCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_add_constant_central_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_add_constant_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_constant_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionAddConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_add_constant_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_add_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionAddConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_add_constant_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_add_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionSetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_set_constant_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_set_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_constant_force[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionSetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_set_constant_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_set_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_constant_torque[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionSetSleepState {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_set_sleep_state[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_set_sleep_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_sleep_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionIsSleeping {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_is_sleeping[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_is_sleeping[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_sleeping")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactCount {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_count[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactLocalPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_local_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_local_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactLocalNormal {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_local_normal[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_local_normal[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_normal")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_impulse[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactLocalShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_local_shape[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_local_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactLocalVelocityAtPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_local_velocity_at_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_local_velocity_at_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_local_velocity_at_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactCollider {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_collider[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_collider[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactColliderPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_collider_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_collider_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactColliderId {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_collider_id[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_collider_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactColliderObject {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_collider_object[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_collider_object[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_object")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactColliderShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_collider_shape[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_collider_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetContactColliderVelocityAtPosition {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_contact_collider_velocity_at_position[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_contact_collider_velocity_at_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contact_collider_velocity_at_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetStep {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_step[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_step[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_step")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionIntegrateForces {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_integrate_forces[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_integrate_forces[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_integrate_forces")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectBodyState3DExtensionGetSpaceState {{
		// HACK: force function generation
		if false { unsafe { physicsdirectbodystate3dextension_gd_get_space_state[T](nil, nil, nil) } }

		func := physicsdirectbodystate3dextension_gd_get_space_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_space_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState2DExtensionIntersectRay {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate2dextension_gd_intersect_ray[T](nil, nil, nil) } }

		func := physicsdirectspacestate2dextension_gd_intersect_ray[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_intersect_ray")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState2DExtensionIntersectPoint {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate2dextension_gd_intersect_point[T](nil, nil, nil) } }

		func := physicsdirectspacestate2dextension_gd_intersect_point[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_intersect_point")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState2DExtensionIntersectShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate2dextension_gd_intersect_shape[T](nil, nil, nil) } }

		func := physicsdirectspacestate2dextension_gd_intersect_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_intersect_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState2DExtensionCastMotion {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate2dextension_gd_cast_motion[T](nil, nil, nil) } }

		func := physicsdirectspacestate2dextension_gd_cast_motion[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cast_motion")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState2DExtensionCollideShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate2dextension_gd_collide_shape[T](nil, nil, nil) } }

		func := physicsdirectspacestate2dextension_gd_collide_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_collide_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState2DExtensionRestInfo {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate2dextension_gd_rest_info[T](nil, nil, nil) } }

		func := physicsdirectspacestate2dextension_gd_rest_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_rest_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState3DExtensionIntersectRay {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate3dextension_gd_intersect_ray[T](nil, nil, nil) } }

		func := physicsdirectspacestate3dextension_gd_intersect_ray[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_intersect_ray")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState3DExtensionIntersectPoint {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate3dextension_gd_intersect_point[T](nil, nil, nil) } }

		func := physicsdirectspacestate3dextension_gd_intersect_point[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_intersect_point")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState3DExtensionIntersectShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate3dextension_gd_intersect_shape[T](nil, nil, nil) } }

		func := physicsdirectspacestate3dextension_gd_intersect_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_intersect_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState3DExtensionCastMotion {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate3dextension_gd_cast_motion[T](nil, nil, nil) } }

		func := physicsdirectspacestate3dextension_gd_cast_motion[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cast_motion")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState3DExtensionCollideShape {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate3dextension_gd_collide_shape[T](nil, nil, nil) } }

		func := physicsdirectspacestate3dextension_gd_collide_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_collide_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState3DExtensionRestInfo {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate3dextension_gd_rest_info[T](nil, nil, nil) } }

		func := physicsdirectspacestate3dextension_gd_rest_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_rest_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsDirectSpaceState3DExtensionGetClosestPointToObjectVolume {{
		// HACK: force function generation
		if false { unsafe { physicsdirectspacestate3dextension_gd_get_closest_point_to_object_volume[T](nil, nil, nil) } }

		func := physicsdirectspacestate3dextension_gd_get_closest_point_to_object_volume[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_closest_point_to_object_volume")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionWorldBoundaryShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_world_boundary_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_world_boundary_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_world_boundary_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSeparationRayShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_separation_ray_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_separation_ray_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_separation_ray_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSegmentShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_segment_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_segment_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_segment_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionCircleShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_circle_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_circle_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_circle_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionRectangleShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_rectangle_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_rectangle_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_rectangle_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionCapsuleShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_capsule_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_capsule_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_capsule_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionConvexPolygonShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_convex_polygon_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_convex_polygon_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_convex_polygon_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionConcavePolygonShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_concave_polygon_shape_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_concave_polygon_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_concave_polygon_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionShapeSetData {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_shape_set_data[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_shape_set_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_set_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionShapeSetCustomSolverBias {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_shape_set_custom_solver_bias[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_shape_set_custom_solver_bias[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_set_custom_solver_bias")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionShapeGetType {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_shape_get_type[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_shape_get_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_get_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionShapeGetData {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_shape_get_data[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_shape_get_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_get_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionShapeGetCustomSolverBias {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_shape_get_custom_solver_bias[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_shape_get_custom_solver_bias[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_get_custom_solver_bias")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionShapeCollide {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_shape_collide[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_shape_collide[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_collide")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceSetActive {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_set_active[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_set_active[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_set_active")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceIsActive {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_is_active[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_is_active[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_is_active")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_set_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_get_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceGetDirectState {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_get_direct_state[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_get_direct_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_direct_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceSetDebugContacts {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_set_debug_contacts[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_set_debug_contacts[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_set_debug_contacts")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceGetContacts {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_get_contacts[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_get_contacts[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_contacts")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSpaceGetContactCount {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_space_get_contact_count[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_space_get_contact_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_contact_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_space[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_space[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaAddShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_add_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_add_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_add_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_shape_transform[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetShapeDisabled {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_shape_disabled[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_shape_disabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_shape_disabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetShapeCount {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_shape_count[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_shape_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_shape_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_shape_transform[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaRemoveShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_remove_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_remove_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_remove_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaClearShapes {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_clear_shapes[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_clear_shapes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_clear_shapes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaAttachObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_attach_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_attach_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_attach_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaAttachCanvasInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_attach_canvas_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_attach_canvas_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_attach_canvas_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetCanvasInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_canvas_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_canvas_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_canvas_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_transform[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_transform[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_collision_layer[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_collision_layer[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_collision_mask[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaGetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_get_collision_mask[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_get_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetMonitorable {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_monitorable[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_monitorable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_monitorable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetPickable {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_pickable[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_pickable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_pickable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetMonitorCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_monitor_callback[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_monitor_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_monitor_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionAreaSetAreaMonitorCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_area_set_area_monitor_callback[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_area_set_area_monitor_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_area_monitor_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_space[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_space[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetMode {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_mode[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetMode {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_mode[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyAddShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_add_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_add_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_shape_transform[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetShapeCount {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_shape_count[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_shape_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_shape_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_shape_transform[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetShapeDisabled {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_shape_disabled[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_shape_disabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_shape_disabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetShapeAsOneWayCollision {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_shape_as_one_way_collision[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_shape_as_one_way_collision[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_shape_as_one_way_collision")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyRemoveShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_remove_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_remove_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_remove_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyClearShapes {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_clear_shapes[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_clear_shapes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_clear_shapes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyAttachObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_attach_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_attach_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_attach_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyAttachCanvasInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_attach_canvas_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_attach_canvas_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_attach_canvas_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetCanvasInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_canvas_instance_id[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_canvas_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_canvas_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetContinuousCollisionDetectionMode {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_continuous_collision_detection_mode[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_continuous_collision_detection_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_continuous_collision_detection_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetContinuousCollisionDetectionMode {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_continuous_collision_detection_mode[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_continuous_collision_detection_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_continuous_collision_detection_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_collision_layer[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_collision_layer[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_collision_mask[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_collision_mask[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetCollisionPriority {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_collision_priority[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_collision_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_collision_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetCollisionPriority {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_collision_priority[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_collision_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyResetMassProperties {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_reset_mass_properties[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_reset_mass_properties[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_reset_mass_properties")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetState {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_state[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetState {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_state[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyApplyCentralImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_apply_central_impulse[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_apply_central_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_central_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyApplyTorqueImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_apply_torque_impulse[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_apply_torque_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_torque_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyApplyImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_apply_impulse[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_apply_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyApplyCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_apply_central_force[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_apply_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyApplyForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_apply_force[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_apply_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyApplyTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_apply_torque[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_apply_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyAddConstantCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_add_constant_central_force[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_add_constant_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_constant_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyAddConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_add_constant_force[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_add_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyAddConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_add_constant_torque[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_add_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_constant_force[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_constant_force[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_constant_torque[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_constant_torque[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetAxisVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_axis_velocity[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_axis_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_axis_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyAddCollisionException {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_add_collision_exception[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_add_collision_exception[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_collision_exception")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyRemoveCollisionException {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_remove_collision_exception[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_remove_collision_exception[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_remove_collision_exception")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetCollisionExceptions {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_collision_exceptions[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_collision_exceptions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_exceptions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetMaxContactsReported {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_max_contacts_reported[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_max_contacts_reported[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_max_contacts_reported")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetMaxContactsReported {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_max_contacts_reported[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_max_contacts_reported[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_max_contacts_reported")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetContactsReportedDepthThreshold {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_contacts_reported_depth_threshold[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_contacts_reported_depth_threshold[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_contacts_reported_depth_threshold")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetContactsReportedDepthThreshold {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_contacts_reported_depth_threshold[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_contacts_reported_depth_threshold[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_contacts_reported_depth_threshold")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetOmitForceIntegration {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_omit_force_integration[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_omit_force_integration[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_omit_force_integration")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyIsOmittingForceIntegration {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_is_omitting_force_integration[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_is_omitting_force_integration[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_is_omitting_force_integration")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetStateSyncCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_state_sync_callback[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_state_sync_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_state_sync_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetForceIntegrationCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_force_integration_callback[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_force_integration_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_force_integration_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyCollideShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_collide_shape[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_collide_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_collide_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodySetPickable {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_set_pickable[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_set_pickable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_pickable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyGetDirectState {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_get_direct_state[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_get_direct_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_direct_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionBodyTestMotion {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_body_test_motion[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_body_test_motion[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_test_motion")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_create[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointClear {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_clear[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_clear[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_clear")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointDisableCollisionsBetweenBodies {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_disable_collisions_between_bodies[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_disable_collisions_between_bodies[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_disable_collisions_between_bodies")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointIsDisabledCollisionsBetweenBodies {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_is_disabled_collisions_between_bodies[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_is_disabled_collisions_between_bodies[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_is_disabled_collisions_between_bodies")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointMakePin {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_make_pin[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_make_pin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_pin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointMakeGroove {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_make_groove[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_make_groove[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_groove")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointMakeDampedSpring {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_make_damped_spring[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_make_damped_spring[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_damped_spring")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionPinJointSetFlag {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_pin_joint_set_flag[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_pin_joint_set_flag[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_set_flag")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionPinJointGetFlag {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_pin_joint_get_flag[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_pin_joint_get_flag[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_get_flag")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionPinJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_pin_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_pin_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionPinJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_pin_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_pin_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionDampedSpringJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_damped_spring_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_damped_spring_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_damped_spring_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionDampedSpringJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_damped_spring_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_damped_spring_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_damped_spring_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionJointGetType {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_joint_get_type[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_joint_get_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_get_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionFreeRid {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_free_rid[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_free_rid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_free_rid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSetActive {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_set_active[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_set_active[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_active")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionInit {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_init[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_init[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_init")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionStep {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_step[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_step[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_step")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionSync {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_sync[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_sync[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_sync")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionFlushQueries {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_flush_queries[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_flush_queries[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_flush_queries")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionEndSync {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_end_sync[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_end_sync[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_end_sync")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionFinish {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_finish[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_finish[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_finish")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionIsFlushingQueries {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_is_flushing_queries[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_is_flushing_queries[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_flushing_queries")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer2DExtensionGetProcessInfo {{
		// HACK: force function generation
		if false { unsafe { physicsserver2dextension_gd_get_process_info[T](nil, nil, nil) } }

		func := physicsserver2dextension_gd_get_process_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_process_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionWorldBoundaryShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_world_boundary_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_world_boundary_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_world_boundary_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSeparationRayShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_separation_ray_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_separation_ray_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_separation_ray_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSphereShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_sphere_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_sphere_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_sphere_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBoxShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_box_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_box_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_box_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionCapsuleShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_capsule_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_capsule_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_capsule_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionCylinderShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_cylinder_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_cylinder_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cylinder_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionConvexPolygonShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_convex_polygon_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_convex_polygon_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_convex_polygon_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionConcavePolygonShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_concave_polygon_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_concave_polygon_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_concave_polygon_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionHeightmapShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_heightmap_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_heightmap_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_heightmap_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionCustomShapeCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_custom_shape_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_custom_shape_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_custom_shape_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionShapeSetData {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_shape_set_data[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_shape_set_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_set_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionShapeSetCustomSolverBias {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_shape_set_custom_solver_bias[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_shape_set_custom_solver_bias[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_set_custom_solver_bias")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionShapeSetMargin {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_shape_set_margin[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_shape_set_margin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_set_margin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionShapeGetMargin {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_shape_get_margin[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_shape_get_margin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_get_margin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionShapeGetType {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_shape_get_type[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_shape_get_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_get_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionShapeGetData {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_shape_get_data[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_shape_get_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_get_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionShapeGetCustomSolverBias {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_shape_get_custom_solver_bias[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_shape_get_custom_solver_bias[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shape_get_custom_solver_bias")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceSetActive {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_set_active[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_set_active[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_set_active")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceIsActive {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_is_active[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_is_active[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_is_active")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceGetDirectState {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_get_direct_state[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_get_direct_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_direct_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceSetDebugContacts {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_set_debug_contacts[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_set_debug_contacts[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_set_debug_contacts")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceGetContacts {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_get_contacts[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_get_contacts[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_contacts")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSpaceGetContactCount {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_space_get_contact_count[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_space_get_contact_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_space_get_contact_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_space[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_space[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaAddShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_add_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_add_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_add_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_shape_transform[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetShapeDisabled {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_shape_disabled[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_shape_disabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_shape_disabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetShapeCount {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_shape_count[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_shape_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_shape_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_shape_transform[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaRemoveShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_remove_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_remove_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_remove_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaClearShapes {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_clear_shapes[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_clear_shapes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_clear_shapes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaAttachObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_attach_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_attach_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_attach_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_transform[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_transform[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_collision_layer[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_collision_layer[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_collision_mask[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaGetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_get_collision_mask[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_get_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_get_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetMonitorable {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_monitorable[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_monitorable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_monitorable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetRayPickable {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_ray_pickable[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_ray_pickable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_ray_pickable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetMonitorCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_monitor_callback[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_monitor_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_monitor_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionAreaSetAreaMonitorCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_area_set_area_monitor_callback[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_area_set_area_monitor_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_area_set_area_monitor_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_space[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_space[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetMode {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_mode[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetMode {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_mode[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyAddShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_add_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_add_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_shape_transform[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetShapeDisabled {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_shape_disabled[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_shape_disabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_shape_disabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetShapeCount {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_shape_count[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_shape_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_shape_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetShapeTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_shape_transform[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_shape_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_shape_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyRemoveShape {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_remove_shape[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_remove_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_remove_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyClearShapes {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_clear_shapes[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_clear_shapes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_clear_shapes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyAttachObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_attach_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_attach_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_attach_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetObjectInstanceId {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_object_instance_id[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_object_instance_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_object_instance_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetEnableContinuousCollisionDetection {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_enable_continuous_collision_detection[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_enable_continuous_collision_detection[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_enable_continuous_collision_detection")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyIsContinuousCollisionDetectionEnabled {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_is_continuous_collision_detection_enabled[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_is_continuous_collision_detection_enabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_is_continuous_collision_detection_enabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_collision_layer[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_collision_layer[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_collision_mask[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_collision_mask[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetCollisionPriority {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_collision_priority[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_collision_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_collision_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetCollisionPriority {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_collision_priority[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_collision_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetUserFlags {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_user_flags[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_user_flags[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_user_flags")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetUserFlags {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_user_flags[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_user_flags[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_user_flags")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyResetMassProperties {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_reset_mass_properties[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_reset_mass_properties[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_reset_mass_properties")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetState {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_state[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetState {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_state[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyApplyCentralImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_apply_central_impulse[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_apply_central_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_central_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyApplyImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_apply_impulse[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_apply_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyApplyTorqueImpulse {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_apply_torque_impulse[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_apply_torque_impulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_torque_impulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyApplyCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_apply_central_force[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_apply_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyApplyForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_apply_force[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_apply_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyApplyTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_apply_torque[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_apply_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_apply_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyAddConstantCentralForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_add_constant_central_force[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_add_constant_central_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_constant_central_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyAddConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_add_constant_force[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_add_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyAddConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_add_constant_torque[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_add_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_constant_force[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetConstantForce {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_constant_force[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_constant_force[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_constant_force")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_constant_torque[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetConstantTorque {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_constant_torque[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_constant_torque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_constant_torque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetAxisVelocity {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_axis_velocity[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_axis_velocity[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_axis_velocity")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetAxisLock {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_axis_lock[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_axis_lock[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_axis_lock")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyIsAxisLocked {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_is_axis_locked[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_is_axis_locked[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_is_axis_locked")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyAddCollisionException {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_add_collision_exception[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_add_collision_exception[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_add_collision_exception")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyRemoveCollisionException {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_remove_collision_exception[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_remove_collision_exception[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_remove_collision_exception")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetCollisionExceptions {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_collision_exceptions[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_collision_exceptions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_collision_exceptions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetMaxContactsReported {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_max_contacts_reported[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_max_contacts_reported[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_max_contacts_reported")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetMaxContactsReported {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_max_contacts_reported[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_max_contacts_reported[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_max_contacts_reported")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetContactsReportedDepthThreshold {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_contacts_reported_depth_threshold[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_contacts_reported_depth_threshold[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_contacts_reported_depth_threshold")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetContactsReportedDepthThreshold {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_contacts_reported_depth_threshold[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_contacts_reported_depth_threshold[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_contacts_reported_depth_threshold")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetOmitForceIntegration {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_omit_force_integration[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_omit_force_integration[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_omit_force_integration")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyIsOmittingForceIntegration {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_is_omitting_force_integration[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_is_omitting_force_integration[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_is_omitting_force_integration")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetStateSyncCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_state_sync_callback[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_state_sync_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_state_sync_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetForceIntegrationCallback {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_force_integration_callback[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_force_integration_callback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_force_integration_callback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodySetRayPickable {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_set_ray_pickable[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_set_ray_pickable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_set_ray_pickable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyTestMotion {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_test_motion[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_test_motion[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_test_motion")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionBodyGetDirectState {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_body_get_direct_state[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_body_get_direct_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_body_get_direct_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyUpdateRenderingServer {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_update_rendering_server[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_update_rendering_server[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_update_rendering_server")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_space[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetSpace {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_space[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_space[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_space")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetRayPickable {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_ray_pickable[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_ray_pickable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_ray_pickable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_collision_layer[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetCollisionLayer {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_collision_layer[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_collision_layer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_collision_layer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_collision_mask[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetCollisionMask {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_collision_mask[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_collision_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_collision_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyAddCollisionException {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_add_collision_exception[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_add_collision_exception[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_add_collision_exception")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyRemoveCollisionException {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_remove_collision_exception[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_remove_collision_exception[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_remove_collision_exception")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetCollisionExceptions {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_collision_exceptions[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_collision_exceptions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_collision_exceptions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetState {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_state[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetState {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_state[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetTransform {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_transform[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetSimulationPrecision {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_simulation_precision[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_simulation_precision[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_simulation_precision")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetSimulationPrecision {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_simulation_precision[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_simulation_precision[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_simulation_precision")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetTotalMass {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_total_mass[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_total_mass[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_total_mass")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetTotalMass {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_total_mass[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_total_mass[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_total_mass")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetLinearStiffness {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_linear_stiffness[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_linear_stiffness[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_linear_stiffness")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetLinearStiffness {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_linear_stiffness[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_linear_stiffness[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_linear_stiffness")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetPressureCoefficient {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_pressure_coefficient[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_pressure_coefficient[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_pressure_coefficient")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetPressureCoefficient {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_pressure_coefficient[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_pressure_coefficient[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_pressure_coefficient")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetDampingCoefficient {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_damping_coefficient[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_damping_coefficient[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_damping_coefficient")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetDampingCoefficient {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_damping_coefficient[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_damping_coefficient[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_damping_coefficient")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetDragCoefficient {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_drag_coefficient[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_drag_coefficient[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_drag_coefficient")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetDragCoefficient {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_drag_coefficient[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_drag_coefficient[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_drag_coefficient")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodySetMesh {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_set_mesh[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_set_mesh[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_set_mesh")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetBounds {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_bounds[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_bounds[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_bounds")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyMovePoint {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_move_point[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_move_point[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_move_point")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyGetPointGlobalPosition {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_get_point_global_position[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_get_point_global_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_get_point_global_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyRemoveAllPinnedPoints {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_remove_all_pinned_points[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_remove_all_pinned_points[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_remove_all_pinned_points")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyPinPoint {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_pin_point[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_pin_point[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_pin_point")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSoftBodyIsPointPinned {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_soft_body_is_point_pinned[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_soft_body_is_point_pinned[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_soft_body_is_point_pinned")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointCreate {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_create[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointClear {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_clear[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_clear[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_clear")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointMakePin {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_make_pin[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_make_pin[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_pin")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionPinJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_pin_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_pin_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionPinJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_pin_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_pin_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionPinJointSetLocalA {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_pin_joint_set_local_a[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_pin_joint_set_local_a[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_set_local_a")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionPinJointGetLocalA {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_pin_joint_get_local_a[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_pin_joint_get_local_a[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_get_local_a")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionPinJointSetLocalB {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_pin_joint_set_local_b[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_pin_joint_set_local_b[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_set_local_b")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionPinJointGetLocalB {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_pin_joint_get_local_b[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_pin_joint_get_local_b[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pin_joint_get_local_b")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointMakeHinge {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_make_hinge[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_make_hinge[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_hinge")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointMakeHingeSimple {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_make_hinge_simple[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_make_hinge_simple[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_hinge_simple")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionHingeJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_hinge_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_hinge_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_hinge_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionHingeJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_hinge_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_hinge_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_hinge_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionHingeJointSetFlag {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_hinge_joint_set_flag[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_hinge_joint_set_flag[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_hinge_joint_set_flag")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionHingeJointGetFlag {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_hinge_joint_get_flag[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_hinge_joint_get_flag[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_hinge_joint_get_flag")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointMakeSlider {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_make_slider[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_make_slider[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_slider")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSliderJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_slider_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_slider_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_slider_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSliderJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_slider_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_slider_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_slider_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointMakeConeTwist {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_make_cone_twist[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_make_cone_twist[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_cone_twist")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionConeTwistJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_cone_twist_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_cone_twist_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cone_twist_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionConeTwistJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_cone_twist_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_cone_twist_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cone_twist_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointMakeGeneric6dof {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_make_generic_6dof[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_make_generic_6dof[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_make_generic_6dof")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionGeneric6dofJointSetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_generic_6dof_joint_set_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_generic_6dof_joint_set_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generic_6dof_joint_set_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionGeneric6dofJointGetParam {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_generic_6dof_joint_get_param[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_generic_6dof_joint_get_param[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generic_6dof_joint_get_param")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionGeneric6dofJointSetFlag {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_generic_6dof_joint_set_flag[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_generic_6dof_joint_set_flag[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generic_6dof_joint_set_flag")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionGeneric6dofJointGetFlag {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_generic_6dof_joint_get_flag[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_generic_6dof_joint_get_flag[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_generic_6dof_joint_get_flag")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointGetType {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_get_type[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_get_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_get_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointSetSolverPriority {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_set_solver_priority[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_set_solver_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_set_solver_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointGetSolverPriority {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_get_solver_priority[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_get_solver_priority[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_get_solver_priority")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointDisableCollisionsBetweenBodies {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_disable_collisions_between_bodies[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_disable_collisions_between_bodies[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_disable_collisions_between_bodies")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionJointIsDisabledCollisionsBetweenBodies {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_joint_is_disabled_collisions_between_bodies[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_joint_is_disabled_collisions_between_bodies[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_joint_is_disabled_collisions_between_bodies")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionFreeRid {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_free_rid[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_free_rid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_free_rid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSetActive {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_set_active[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_set_active[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_active")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionInit {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_init[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_init[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_init")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionStep {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_step[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_step[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_step")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionSync {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_sync[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_sync[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_sync")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionFlushQueries {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_flush_queries[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_flush_queries[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_flush_queries")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionEndSync {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_end_sync[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_end_sync[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_end_sync")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionFinish {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_finish[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_finish[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_finish")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionIsFlushingQueries {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_is_flushing_queries[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_is_flushing_queries[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_flushing_queries")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DExtensionGetProcessInfo {{
		// HACK: force function generation
		if false { unsafe { physicsserver3dextension_gd_get_process_info[T](nil, nil, nil) } }

		func := physicsserver3dextension_gd_get_process_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_process_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DRenderingServerHandlerSetVertex {{
		// HACK: force function generation
		if false { unsafe { physicsserver3drenderingserverhandler_gd_set_vertex[T](nil, nil, nil) } }

		func := physicsserver3drenderingserverhandler_gd_set_vertex[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_vertex")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DRenderingServerHandlerSetNormal {{
		// HACK: force function generation
		if false { unsafe { physicsserver3drenderingserverhandler_gd_set_normal[T](nil, nil, nil) } }

		func := physicsserver3drenderingserverhandler_gd_set_normal[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_normal")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPhysicsServer3DRenderingServerHandlerSetAabb {{
		// HACK: force function generation
		if false { unsafe { physicsserver3drenderingserverhandler_gd_set_aabb[T](nil, nil, nil) } }

		func := physicsserver3drenderingserverhandler_gd_set_aabb[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_aabb")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IPrimitiveMeshCreateMeshArray {{
		// HACK: force function generation
		if false { unsafe { primitivemesh_gd_create_mesh_array[T](nil, nil, nil) } }

		func := primitivemesh_gd_create_mesh_array[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_mesh_array")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRangeValueChanged {{
		// HACK: force function generation
		if false { unsafe { range_gd_value_changed[T](nil, nil, nil) } }

		func := range_gd_value_changed[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_value_changed")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderDataExtensionGetRenderSceneBuffers {{
		// HACK: force function generation
		if false { unsafe { renderdataextension_gd_get_render_scene_buffers[T](nil, nil, nil) } }

		func := renderdataextension_gd_get_render_scene_buffers[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_render_scene_buffers")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderDataExtensionGetRenderSceneData {{
		// HACK: force function generation
		if false { unsafe { renderdataextension_gd_get_render_scene_data[T](nil, nil, nil) } }

		func := renderdataextension_gd_get_render_scene_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_render_scene_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderDataExtensionGetEnvironment {{
		// HACK: force function generation
		if false { unsafe { renderdataextension_gd_get_environment[T](nil, nil, nil) } }

		func := renderdataextension_gd_get_environment[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_environment")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderDataExtensionGetCameraAttributes {{
		// HACK: force function generation
		if false { unsafe { renderdataextension_gd_get_camera_attributes[T](nil, nil, nil) } }

		func := renderdataextension_gd_get_camera_attributes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_camera_attributes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneBuffersExtensionConfigure {{
		// HACK: force function generation
		if false { unsafe { renderscenebuffersextension_gd_configure[T](nil, nil, nil) } }

		func := renderscenebuffersextension_gd_configure[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_configure")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneBuffersExtensionSetFsrSharpness {{
		// HACK: force function generation
		if false { unsafe { renderscenebuffersextension_gd_set_fsr_sharpness[T](nil, nil, nil) } }

		func := renderscenebuffersextension_gd_set_fsr_sharpness[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_fsr_sharpness")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneBuffersExtensionSetTextureMipmapBias {{
		// HACK: force function generation
		if false { unsafe { renderscenebuffersextension_gd_set_texture_mipmap_bias[T](nil, nil, nil) } }

		func := renderscenebuffersextension_gd_set_texture_mipmap_bias[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_texture_mipmap_bias")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneBuffersExtensionSetAnisotropicFilteringLevel {{
		// HACK: force function generation
		if false { unsafe { renderscenebuffersextension_gd_set_anisotropic_filtering_level[T](nil, nil, nil) } }

		func := renderscenebuffersextension_gd_set_anisotropic_filtering_level[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_anisotropic_filtering_level")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneBuffersExtensionSetUseDebanding {{
		// HACK: force function generation
		if false { unsafe { renderscenebuffersextension_gd_set_use_debanding[T](nil, nil, nil) } }

		func := renderscenebuffersextension_gd_set_use_debanding[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_use_debanding")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneDataExtensionGetCamTransform {{
		// HACK: force function generation
		if false { unsafe { renderscenedataextension_gd_get_cam_transform[T](nil, nil, nil) } }

		func := renderscenedataextension_gd_get_cam_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_cam_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneDataExtensionGetCamProjection {{
		// HACK: force function generation
		if false { unsafe { renderscenedataextension_gd_get_cam_projection[T](nil, nil, nil) } }

		func := renderscenedataextension_gd_get_cam_projection[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_cam_projection")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneDataExtensionGetViewCount {{
		// HACK: force function generation
		if false { unsafe { renderscenedataextension_gd_get_view_count[T](nil, nil, nil) } }

		func := renderscenedataextension_gd_get_view_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_view_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneDataExtensionGetViewEyeOffset {{
		// HACK: force function generation
		if false { unsafe { renderscenedataextension_gd_get_view_eye_offset[T](nil, nil, nil) } }

		func := renderscenedataextension_gd_get_view_eye_offset[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_view_eye_offset")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneDataExtensionGetViewProjection {{
		// HACK: force function generation
		if false { unsafe { renderscenedataextension_gd_get_view_projection[T](nil, nil, nil) } }

		func := renderscenedataextension_gd_get_view_projection[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_view_projection")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRenderSceneDataExtensionGetUniformBuffer {{
		// HACK: force function generation
		if false { unsafe { renderscenedataextension_gd_get_uniform_buffer[T](nil, nil, nil) } }

		func := renderscenedataextension_gd_get_uniform_buffer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_uniform_buffer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceSetupLocalToScene {{
		// HACK: force function generation
		if false { unsafe { resource_gd_setup_local_to_scene[T](nil, nil, nil) } }

		func := resource_gd_setup_local_to_scene[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_setup_local_to_scene")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceGetRid {{
		// HACK: force function generation
		if false { unsafe { resource_gd_get_rid[T](nil, nil, nil) } }

		func := resource_gd_get_rid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_rid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceResetState {{
		// HACK: force function generation
		if false { unsafe { resource_gd_reset_state[T](nil, nil, nil) } }

		func := resource_gd_reset_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_reset_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceSetPathCache {{
		// HACK: force function generation
		if false { unsafe { resource_gd_set_path_cache[T](nil, nil, nil) } }

		func := resource_gd_set_path_cache[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_path_cache")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderGetRecognizedExtensions {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_get_recognized_extensions[T](nil, nil, nil) } }

		func := resourceformatloader_gd_get_recognized_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_recognized_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderRecognizePath {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_recognize_path[T](nil, nil, nil) } }

		func := resourceformatloader_gd_recognize_path[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_recognize_path")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderHandlesType {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_handles_type[T](nil, nil, nil) } }

		func := resourceformatloader_gd_handles_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handles_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderGetResourceType {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_get_resource_type[T](nil, nil, nil) } }

		func := resourceformatloader_gd_get_resource_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_resource_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderGetResourceScriptClass {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_get_resource_script_class[T](nil, nil, nil) } }

		func := resourceformatloader_gd_get_resource_script_class[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_resource_script_class")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderGetResourceUid {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_get_resource_uid[T](nil, nil, nil) } }

		func := resourceformatloader_gd_get_resource_uid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_resource_uid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderGetDependencies {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_get_dependencies[T](nil, nil, nil) } }

		func := resourceformatloader_gd_get_dependencies[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_dependencies")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderRenameDependencies {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_rename_dependencies[T](nil, nil, nil) } }

		func := resourceformatloader_gd_rename_dependencies[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_rename_dependencies")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderExists {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_exists[T](nil, nil, nil) } }

		func := resourceformatloader_gd_exists[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_exists")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderGetClassesUsed {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_get_classes_used[T](nil, nil, nil) } }

		func := resourceformatloader_gd_get_classes_used[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_classes_used")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatLoaderLoad {{
		// HACK: force function generation
		if false { unsafe { resourceformatloader_gd_load[T](nil, nil, nil) } }

		func := resourceformatloader_gd_load[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_load")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatSaverSave {{
		// HACK: force function generation
		if false { unsafe { resourceformatsaver_gd_save[T](nil, nil, nil) } }

		func := resourceformatsaver_gd_save[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_save")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatSaverSetUid {{
		// HACK: force function generation
		if false { unsafe { resourceformatsaver_gd_set_uid[T](nil, nil, nil) } }

		func := resourceformatsaver_gd_set_uid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_uid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatSaverRecognize {{
		// HACK: force function generation
		if false { unsafe { resourceformatsaver_gd_recognize[T](nil, nil, nil) } }

		func := resourceformatsaver_gd_recognize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_recognize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatSaverGetRecognizedExtensions {{
		// HACK: force function generation
		if false { unsafe { resourceformatsaver_gd_get_recognized_extensions[T](nil, nil, nil) } }

		func := resourceformatsaver_gd_get_recognized_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_recognized_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IResourceFormatSaverRecognizePath {{
		// HACK: force function generation
		if false { unsafe { resourceformatsaver_gd_recognize_path[T](nil, nil, nil) } }

		func := resourceformatsaver_gd_recognize_path[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_recognize_path")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRichTextEffectProcessCustomFx {{
		// HACK: force function generation
		if false { unsafe { richtexteffect_gd_process_custom_fx[T](nil, nil, nil) } }

		func := richtexteffect_gd_process_custom_fx[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process_custom_fx")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRigidBody2DIntegrateForces {{
		// HACK: force function generation
		if false { unsafe { rigidbody2d_gd_integrate_forces[T](nil, nil, nil) } }

		func := rigidbody2d_gd_integrate_forces[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_integrate_forces")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IRigidBody3DIntegrateForces {{
		// HACK: force function generation
		if false { unsafe { rigidbody3d_gd_integrate_forces[T](nil, nil, nil) } }

		func := rigidbody3d_gd_integrate_forces[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_integrate_forces")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionEditorCanReloadFromFile {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_editor_can_reload_from_file[T](nil, nil, nil) } }

		func := scriptextension_gd_editor_can_reload_from_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_editor_can_reload_from_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionPlaceholderErased {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_placeholder_erased[T](nil, nil, nil) } }

		func := scriptextension_gd_placeholder_erased[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_placeholder_erased")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionCanInstantiate {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_can_instantiate[T](nil, nil, nil) } }

		func := scriptextension_gd_can_instantiate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_instantiate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetBaseScript {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_base_script[T](nil, nil, nil) } }

		func := scriptextension_gd_get_base_script[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_base_script")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetGlobalName {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_global_name[T](nil, nil, nil) } }

		func := scriptextension_gd_get_global_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_global_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionInheritsScript {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_inherits_script[T](nil, nil, nil) } }

		func := scriptextension_gd_inherits_script[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_inherits_script")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetInstanceBaseType {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_instance_base_type[T](nil, nil, nil) } }

		func := scriptextension_gd_get_instance_base_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_instance_base_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionInstanceCreate {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_instance_create[T](nil, nil, nil) } }

		func := scriptextension_gd_instance_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_instance_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionPlaceholderInstanceCreate {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_placeholder_instance_create[T](nil, nil, nil) } }

		func := scriptextension_gd_placeholder_instance_create[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_placeholder_instance_create")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionInstanceHas {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_instance_has[T](nil, nil, nil) } }

		func := scriptextension_gd_instance_has[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_instance_has")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionHasSourceCode {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_has_source_code[T](nil, nil, nil) } }

		func := scriptextension_gd_has_source_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_source_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetSourceCode {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_source_code[T](nil, nil, nil) } }

		func := scriptextension_gd_get_source_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_source_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionSetSourceCode {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_set_source_code[T](nil, nil, nil) } }

		func := scriptextension_gd_set_source_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_source_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionReload {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_reload[T](nil, nil, nil) } }

		func := scriptextension_gd_reload[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_reload")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetDocClassName {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_doc_class_name[T](nil, nil, nil) } }

		func := scriptextension_gd_get_doc_class_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_doc_class_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetDocumentation {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_documentation[T](nil, nil, nil) } }

		func := scriptextension_gd_get_documentation[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_documentation")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetClassIconPath {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_class_icon_path[T](nil, nil, nil) } }

		func := scriptextension_gd_get_class_icon_path[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_class_icon_path")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionHasMethod {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_has_method[T](nil, nil, nil) } }

		func := scriptextension_gd_has_method[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_method")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionHasStaticMethod {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_has_static_method[T](nil, nil, nil) } }

		func := scriptextension_gd_has_static_method[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_static_method")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetScriptMethodArgumentCount {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_script_method_argument_count[T](nil, nil, nil) } }

		func := scriptextension_gd_get_script_method_argument_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_script_method_argument_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetMethodInfo {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_method_info[T](nil, nil, nil) } }

		func := scriptextension_gd_get_method_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_method_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionIsTool {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_is_tool[T](nil, nil, nil) } }

		func := scriptextension_gd_is_tool[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_tool")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionIsValid {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_is_valid[T](nil, nil, nil) } }

		func := scriptextension_gd_is_valid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_valid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionIsAbstract {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_is_abstract[T](nil, nil, nil) } }

		func := scriptextension_gd_is_abstract[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_abstract")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetLanguage {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_language[T](nil, nil, nil) } }

		func := scriptextension_gd_get_language[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_language")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionHasScriptSignal {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_has_script_signal[T](nil, nil, nil) } }

		func := scriptextension_gd_has_script_signal[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_script_signal")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetScriptSignalList {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_script_signal_list[T](nil, nil, nil) } }

		func := scriptextension_gd_get_script_signal_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_script_signal_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionHasPropertyDefaultValue {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_has_property_default_value[T](nil, nil, nil) } }

		func := scriptextension_gd_has_property_default_value[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_property_default_value")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetPropertyDefaultValue {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_property_default_value[T](nil, nil, nil) } }

		func := scriptextension_gd_get_property_default_value[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_property_default_value")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionUpdateExports {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_update_exports[T](nil, nil, nil) } }

		func := scriptextension_gd_update_exports[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_update_exports")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetScriptMethodList {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_script_method_list[T](nil, nil, nil) } }

		func := scriptextension_gd_get_script_method_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_script_method_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetScriptPropertyList {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_script_property_list[T](nil, nil, nil) } }

		func := scriptextension_gd_get_script_property_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_script_property_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetMemberLine {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_member_line[T](nil, nil, nil) } }

		func := scriptextension_gd_get_member_line[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_member_line")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetConstants {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_constants[T](nil, nil, nil) } }

		func := scriptextension_gd_get_constants[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_constants")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetMembers {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_members[T](nil, nil, nil) } }

		func := scriptextension_gd_get_members[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_members")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionIsPlaceholderFallbackEnabled {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_is_placeholder_fallback_enabled[T](nil, nil, nil) } }

		func := scriptextension_gd_is_placeholder_fallback_enabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_placeholder_fallback_enabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptExtensionGetRpcConfig {{
		// HACK: force function generation
		if false { unsafe { scriptextension_gd_get_rpc_config[T](nil, nil, nil) } }

		func := scriptextension_gd_get_rpc_config[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_rpc_config")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetName {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_name[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionInit {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_init[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_init[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_init")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetType {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_type[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetExtension {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_extension[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_extension[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_extension")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionFinish {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_finish[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_finish[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_finish")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetReservedWords {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_reserved_words[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_reserved_words[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_reserved_words")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionIsControlFlowKeyword {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_is_control_flow_keyword[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_is_control_flow_keyword[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_control_flow_keyword")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetCommentDelimiters {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_comment_delimiters[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_comment_delimiters[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_comment_delimiters")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetDocCommentDelimiters {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_doc_comment_delimiters[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_doc_comment_delimiters[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_doc_comment_delimiters")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetStringDelimiters {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_string_delimiters[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_string_delimiters[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_string_delimiters")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionMakeTemplate {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_make_template[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_make_template[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_make_template")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetBuiltInTemplates {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_built_in_templates[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_built_in_templates[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_built_in_templates")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionIsUsingTemplates {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_is_using_templates[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_is_using_templates[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_using_templates")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionValidate {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_validate[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_validate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_validate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionValidatePath {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_validate_path[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_validate_path[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_validate_path")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionCreateScript {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_create_script[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_create_script[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_script")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionHasNamedClasses {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_has_named_classes[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_has_named_classes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_named_classes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionSupportsBuiltinMode {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_supports_builtin_mode[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_supports_builtin_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_supports_builtin_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionSupportsDocumentation {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_supports_documentation[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_supports_documentation[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_supports_documentation")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionCanInheritFromFile {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_can_inherit_from_file[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_can_inherit_from_file[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_inherit_from_file")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionFindFunction {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_find_function[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_find_function[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_find_function")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionMakeFunction {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_make_function[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_make_function[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_make_function")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionCanMakeFunction {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_can_make_function[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_can_make_function[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_can_make_function")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionOpenInExternalEditor {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_open_in_external_editor[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_open_in_external_editor[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_open_in_external_editor")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionOverridesExternalEditor {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_overrides_external_editor[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_overrides_external_editor[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_overrides_external_editor")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionPreferredFileNameCasing {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_preferred_file_name_casing[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_preferred_file_name_casing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_preferred_file_name_casing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionCompleteCode {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_complete_code[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_complete_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_complete_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionLookupCode {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_lookup_code[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_lookup_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_lookup_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionAutoIndentCode {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_auto_indent_code[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_auto_indent_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_auto_indent_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionAddGlobalConstant {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_add_global_constant[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_add_global_constant[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_global_constant")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionAddNamedGlobalConstant {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_add_named_global_constant[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_add_named_global_constant[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_named_global_constant")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionRemoveNamedGlobalConstant {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_remove_named_global_constant[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_remove_named_global_constant[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_remove_named_global_constant")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionThreadEnter {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_thread_enter[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_thread_enter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_thread_enter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionThreadExit {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_thread_exit[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_thread_exit[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_thread_exit")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetError {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_error[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_error[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_error")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetStackLevelCount {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_stack_level_count[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_stack_level_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_stack_level_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetStackLevelLine {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_stack_level_line[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_stack_level_line[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_stack_level_line")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetStackLevelFunction {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_stack_level_function[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_stack_level_function[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_stack_level_function")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetStackLevelSource {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_stack_level_source[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_stack_level_source[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_stack_level_source")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetStackLevelLocals {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_stack_level_locals[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_stack_level_locals[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_stack_level_locals")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetStackLevelMembers {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_stack_level_members[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_stack_level_members[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_stack_level_members")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetStackLevelInstance {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_stack_level_instance[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_stack_level_instance[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_stack_level_instance")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetGlobals {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_globals[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_globals[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_globals")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugParseStackLevelExpression {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_parse_stack_level_expression[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_parse_stack_level_expression[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_parse_stack_level_expression")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionDebugGetCurrentStackInfo {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_debug_get_current_stack_info[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_debug_get_current_stack_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_debug_get_current_stack_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionReloadAllScripts {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_reload_all_scripts[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_reload_all_scripts[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_reload_all_scripts")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionReloadScripts {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_reload_scripts[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_reload_scripts[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_reload_scripts")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionReloadToolScript {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_reload_tool_script[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_reload_tool_script[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_reload_tool_script")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetRecognizedExtensions {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_recognized_extensions[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_recognized_extensions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_recognized_extensions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetPublicFunctions {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_public_functions[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_public_functions[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_public_functions")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetPublicConstants {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_public_constants[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_public_constants[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_public_constants")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetPublicAnnotations {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_public_annotations[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_public_annotations[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_public_annotations")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionProfilingStart {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_profiling_start[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_profiling_start[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_profiling_start")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionProfilingStop {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_profiling_stop[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_profiling_stop[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_profiling_stop")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionProfilingSetSaveNativeCalls {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_profiling_set_save_native_calls[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_profiling_set_save_native_calls[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_profiling_set_save_native_calls")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionProfilingGetAccumulatedData {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_profiling_get_accumulated_data[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_profiling_get_accumulated_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_profiling_get_accumulated_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionProfilingGetFrameData {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_profiling_get_frame_data[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_profiling_get_frame_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_profiling_get_frame_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionFrame {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_frame[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_frame[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_frame")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionHandlesGlobalClassType {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_handles_global_class_type[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_handles_global_class_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handles_global_class_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IScriptLanguageExtensionGetGlobalClassName {{
		// HACK: force function generation
		if false { unsafe { scriptlanguageextension_gd_get_global_class_name[T](nil, nil, nil) } }

		func := scriptlanguageextension_gd_get_global_class_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_global_class_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISkeletonModification2DExecute {{
		// HACK: force function generation
		if false { unsafe { skeletonmodification2d_gd_execute[T](nil, nil, nil) } }

		func := skeletonmodification2d_gd_execute[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_execute")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISkeletonModification2DSetupModification {{
		// HACK: force function generation
		if false { unsafe { skeletonmodification2d_gd_setup_modification[T](nil, nil, nil) } }

		func := skeletonmodification2d_gd_setup_modification[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_setup_modification")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISkeletonModification2DDrawEditorGizmo {{
		// HACK: force function generation
		if false { unsafe { skeletonmodification2d_gd_draw_editor_gizmo[T](nil, nil, nil) } }

		func := skeletonmodification2d_gd_draw_editor_gizmo[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw_editor_gizmo")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISkeletonModifier3DProcessModificationWithDelta {{
		// HACK: force function generation
		if false { unsafe { skeletonmodifier3d_gd_process_modification_with_delta[T](nil, nil, nil) } }

		func := skeletonmodifier3d_gd_process_modification_with_delta[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process_modification_with_delta")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISkeletonModifier3DProcessModification {{
		// HACK: force function generation
		if false { unsafe { skeletonmodifier3d_gd_process_modification[T](nil, nil, nil) } }

		func := skeletonmodifier3d_gd_process_modification[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process_modification")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStreamPeerExtensionGetData {{
		// HACK: force function generation
		if false { unsafe { streampeerextension_gd_get_data[T](nil, nil, nil) } }

		func := streampeerextension_gd_get_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStreamPeerExtensionGetPartialData {{
		// HACK: force function generation
		if false { unsafe { streampeerextension_gd_get_partial_data[T](nil, nil, nil) } }

		func := streampeerextension_gd_get_partial_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_partial_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStreamPeerExtensionPutData {{
		// HACK: force function generation
		if false { unsafe { streampeerextension_gd_put_data[T](nil, nil, nil) } }

		func := streampeerextension_gd_put_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_put_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStreamPeerExtensionPutPartialData {{
		// HACK: force function generation
		if false { unsafe { streampeerextension_gd_put_partial_data[T](nil, nil, nil) } }

		func := streampeerextension_gd_put_partial_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_put_partial_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStreamPeerExtensionGetAvailableBytes {{
		// HACK: force function generation
		if false { unsafe { streampeerextension_gd_get_available_bytes[T](nil, nil, nil) } }

		func := streampeerextension_gd_get_available_bytes[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_available_bytes")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStyleBoxDraw {{
		// HACK: force function generation
		if false { unsafe { stylebox_gd_draw[T](nil, nil, nil) } }

		func := stylebox_gd_draw[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStyleBoxGetDrawRect {{
		// HACK: force function generation
		if false { unsafe { stylebox_gd_get_draw_rect[T](nil, nil, nil) } }

		func := stylebox_gd_get_draw_rect[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_draw_rect")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStyleBoxGetMinimumSize {{
		// HACK: force function generation
		if false { unsafe { stylebox_gd_get_minimum_size[T](nil, nil, nil) } }

		func := stylebox_gd_get_minimum_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_minimum_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IStyleBoxTestMask {{
		// HACK: force function generation
		if false { unsafe { stylebox_gd_test_mask[T](nil, nil, nil) } }

		func := stylebox_gd_test_mask[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_test_mask")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISubViewportContainerPropagateInputEvent {{
		// HACK: force function generation
		if false { unsafe { subviewportcontainer_gd_propagate_input_event[T](nil, nil, nil) } }

		func := subviewportcontainer_gd_propagate_input_event[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_propagate_input_event")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISyntaxHighlighterGetLineSyntaxHighlighting {{
		// HACK: force function generation
		if false { unsafe { syntaxhighlighter_gd_get_line_syntax_highlighting[T](nil, nil, nil) } }

		func := syntaxhighlighter_gd_get_line_syntax_highlighting[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_line_syntax_highlighting")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISyntaxHighlighterClearHighlightingCache {{
		// HACK: force function generation
		if false { unsafe { syntaxhighlighter_gd_clear_highlighting_cache[T](nil, nil, nil) } }

		func := syntaxhighlighter_gd_clear_highlighting_cache[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_clear_highlighting_cache")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ISyntaxHighlighterUpdateCache {{
		// HACK: force function generation
		if false { unsafe { syntaxhighlighter_gd_update_cache[T](nil, nil, nil) } }

		func := syntaxhighlighter_gd_update_cache[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_update_cache")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextEditHandleUnicodeInput {{
		// HACK: force function generation
		if false { unsafe { textedit_gd_handle_unicode_input[T](nil, nil, nil) } }

		func := textedit_gd_handle_unicode_input[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_handle_unicode_input")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextEditBackspace {{
		// HACK: force function generation
		if false { unsafe { textedit_gd_backspace[T](nil, nil, nil) } }

		func := textedit_gd_backspace[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_backspace")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextEditCut {{
		// HACK: force function generation
		if false { unsafe { textedit_gd_cut[T](nil, nil, nil) } }

		func := textedit_gd_cut[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cut")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextEditCopy {{
		// HACK: force function generation
		if false { unsafe { textedit_gd_copy[T](nil, nil, nil) } }

		func := textedit_gd_copy[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_copy")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextEditPaste {{
		// HACK: force function generation
		if false { unsafe { textedit_gd_paste[T](nil, nil, nil) } }

		func := textedit_gd_paste[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_paste")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextEditPastePrimaryClipboard {{
		// HACK: force function generation
		if false { unsafe { textedit_gd_paste_primary_clipboard[T](nil, nil, nil) } }

		func := textedit_gd_paste_primary_clipboard[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_paste_primary_clipboard")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionHasFeature {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_has_feature[T](nil, nil, nil) } }

		func := textserverextension_gd_has_feature[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_feature")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionGetName {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_get_name[T](nil, nil, nil) } }

		func := textserverextension_gd_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionGetFeatures {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_get_features[T](nil, nil, nil) } }

		func := textserverextension_gd_get_features[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_features")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFreeRid {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_free_rid[T](nil, nil, nil) } }

		func := textserverextension_gd_free_rid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_free_rid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionHas {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_has[T](nil, nil, nil) } }

		func := textserverextension_gd_has[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionLoadSupportData {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_load_support_data[T](nil, nil, nil) } }

		func := textserverextension_gd_load_support_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_load_support_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionGetSupportDataFilename {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_get_support_data_filename[T](nil, nil, nil) } }

		func := textserverextension_gd_get_support_data_filename[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_support_data_filename")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionGetSupportDataInfo {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_get_support_data_info[T](nil, nil, nil) } }

		func := textserverextension_gd_get_support_data_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_support_data_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionSaveSupportData {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_save_support_data[T](nil, nil, nil) } }

		func := textserverextension_gd_save_support_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_save_support_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionGetSupportData {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_get_support_data[T](nil, nil, nil) } }

		func := textserverextension_gd_get_support_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_support_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionIsLocaleRightToLeft {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_is_locale_right_to_left[T](nil, nil, nil) } }

		func := textserverextension_gd_is_locale_right_to_left[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_locale_right_to_left")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionNameToTag {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_name_to_tag[T](nil, nil, nil) } }

		func := textserverextension_gd_name_to_tag[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_name_to_tag")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionTagToName {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_tag_to_name[T](nil, nil, nil) } }

		func := textserverextension_gd_tag_to_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_tag_to_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionCreateFont {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_create_font[T](nil, nil, nil) } }

		func := textserverextension_gd_create_font[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_font")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionCreateFontLinkedVariation {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_create_font_linked_variation[T](nil, nil, nil) } }

		func := textserverextension_gd_create_font_linked_variation[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_font_linked_variation")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetData {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_data[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetDataPtr {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_data_ptr[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_data_ptr[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_data_ptr")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetFaceIndex {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_face_index[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_face_index[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_face_index")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetFaceIndex {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_face_index[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_face_index[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_face_index")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetFaceCount {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_face_count[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_face_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_face_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetStyle {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_style[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_style[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_style")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetStyle {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_style[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_style[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_style")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetName {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_name[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetName {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_name[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetOtNameStrings {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_ot_name_strings[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_ot_name_strings[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_ot_name_strings")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetStyleName {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_style_name[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_style_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_style_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetStyleName {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_style_name[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_style_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_style_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetWeight {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_weight[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_weight[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_weight")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetWeight {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_weight[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_weight[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_weight")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetStretch {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_stretch[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_stretch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_stretch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetStretch {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_stretch[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_stretch[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_stretch")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetAntialiasing {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_antialiasing[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_antialiasing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_antialiasing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetAntialiasing {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_antialiasing[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_antialiasing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_antialiasing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetDisableEmbeddedBitmaps {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_disable_embedded_bitmaps[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_disable_embedded_bitmaps[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_disable_embedded_bitmaps")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetDisableEmbeddedBitmaps {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_disable_embedded_bitmaps[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_disable_embedded_bitmaps[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_disable_embedded_bitmaps")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetGenerateMipmaps {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_generate_mipmaps[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_generate_mipmaps[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_generate_mipmaps")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGenerateMipmaps {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_generate_mipmaps[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_generate_mipmaps[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_generate_mipmaps")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetMultichannelSignedDistanceField {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_multichannel_signed_distance_field[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_multichannel_signed_distance_field[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_multichannel_signed_distance_field")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontIsMultichannelSignedDistanceField {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_is_multichannel_signed_distance_field[T](nil, nil, nil) } }

		func := textserverextension_gd_font_is_multichannel_signed_distance_field[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_is_multichannel_signed_distance_field")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetMsdfPixelRange {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_msdf_pixel_range[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_msdf_pixel_range[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_msdf_pixel_range")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetMsdfPixelRange {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_msdf_pixel_range[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_msdf_pixel_range[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_msdf_pixel_range")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetMsdfSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_msdf_size[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_msdf_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_msdf_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetMsdfSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_msdf_size[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_msdf_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_msdf_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetFixedSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_fixed_size[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_fixed_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_fixed_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetFixedSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_fixed_size[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_fixed_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_fixed_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetFixedSizeScaleMode {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_fixed_size_scale_mode[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_fixed_size_scale_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_fixed_size_scale_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetFixedSizeScaleMode {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_fixed_size_scale_mode[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_fixed_size_scale_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_fixed_size_scale_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetAllowSystemFallback {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_allow_system_fallback[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_allow_system_fallback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_allow_system_fallback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontIsAllowSystemFallback {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_is_allow_system_fallback[T](nil, nil, nil) } }

		func := textserverextension_gd_font_is_allow_system_fallback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_is_allow_system_fallback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetForceAutohinter {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_force_autohinter[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_force_autohinter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_force_autohinter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontIsForceAutohinter {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_is_force_autohinter[T](nil, nil, nil) } }

		func := textserverextension_gd_font_is_force_autohinter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_is_force_autohinter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetModulateColorGlyphs {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_modulate_color_glyphs[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_modulate_color_glyphs[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_modulate_color_glyphs")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontIsModulateColorGlyphs {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_is_modulate_color_glyphs[T](nil, nil, nil) } }

		func := textserverextension_gd_font_is_modulate_color_glyphs[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_is_modulate_color_glyphs")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetHinting {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_hinting[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_hinting[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_hinting")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetHinting {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_hinting[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_hinting[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_hinting")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetSubpixelPositioning {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_subpixel_positioning[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_subpixel_positioning[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_subpixel_positioning")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetSubpixelPositioning {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_subpixel_positioning[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_subpixel_positioning[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_subpixel_positioning")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetKeepRoundingRemainders {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_keep_rounding_remainders[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_keep_rounding_remainders[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_keep_rounding_remainders")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetKeepRoundingRemainders {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_keep_rounding_remainders[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_keep_rounding_remainders[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_keep_rounding_remainders")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetEmbolden {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_embolden[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_embolden[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_embolden")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetEmbolden {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_embolden[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_embolden[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_embolden")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetSpacing {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_spacing[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_spacing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_spacing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetSpacing {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_spacing[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_spacing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_spacing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetBaselineOffset {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_baseline_offset[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_baseline_offset[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_baseline_offset")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetBaselineOffset {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_baseline_offset[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_baseline_offset[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_baseline_offset")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetTransform {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_transform[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetTransform {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_transform[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetVariationCoordinates {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_variation_coordinates[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_variation_coordinates[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_variation_coordinates")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetVariationCoordinates {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_variation_coordinates[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_variation_coordinates[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_variation_coordinates")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetOversampling {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_oversampling[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_oversampling[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_oversampling")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetOversampling {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_oversampling[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_oversampling[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_oversampling")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetSizeCacheList {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_size_cache_list[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_size_cache_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_size_cache_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontClearSizeCache {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_clear_size_cache[T](nil, nil, nil) } }

		func := textserverextension_gd_font_clear_size_cache[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_clear_size_cache")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRemoveSizeCache {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_remove_size_cache[T](nil, nil, nil) } }

		func := textserverextension_gd_font_remove_size_cache[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_remove_size_cache")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetAscent {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_ascent[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_ascent[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_ascent")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetAscent {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_ascent[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_ascent[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_ascent")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetDescent {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_descent[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_descent[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_descent")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetDescent {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_descent[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_descent[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_descent")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetUnderlinePosition {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_underline_position[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_underline_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_underline_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetUnderlinePosition {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_underline_position[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_underline_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_underline_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetUnderlineThickness {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_underline_thickness[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_underline_thickness[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_underline_thickness")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetUnderlineThickness {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_underline_thickness[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_underline_thickness[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_underline_thickness")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetScale {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_scale[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_scale[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_scale")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetScale {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_scale[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_scale[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_scale")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetTextureCount {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_texture_count[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_texture_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_texture_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontClearTextures {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_clear_textures[T](nil, nil, nil) } }

		func := textserverextension_gd_font_clear_textures[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_clear_textures")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRemoveTexture {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_remove_texture[T](nil, nil, nil) } }

		func := textserverextension_gd_font_remove_texture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_remove_texture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetTextureImage {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_texture_image[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_texture_image[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_texture_image")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetTextureImage {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_texture_image[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_texture_image[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_texture_image")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetTextureOffsets {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_texture_offsets[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_texture_offsets[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_texture_offsets")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetTextureOffsets {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_texture_offsets[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_texture_offsets[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_texture_offsets")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphList {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_list[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontClearGlyphs {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_clear_glyphs[T](nil, nil, nil) } }

		func := textserverextension_gd_font_clear_glyphs[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_clear_glyphs")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRemoveGlyph {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_remove_glyph[T](nil, nil, nil) } }

		func := textserverextension_gd_font_remove_glyph[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_remove_glyph")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphAdvance {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_advance[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_advance[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_advance")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetGlyphAdvance {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_glyph_advance[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_glyph_advance[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_glyph_advance")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphOffset {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_offset[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_offset[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_offset")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetGlyphOffset {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_glyph_offset[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_glyph_offset[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_glyph_offset")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_size[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetGlyphSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_glyph_size[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_glyph_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_glyph_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphUvRect {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_uv_rect[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_uv_rect[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_uv_rect")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetGlyphUvRect {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_glyph_uv_rect[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_glyph_uv_rect[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_glyph_uv_rect")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphTextureIdx {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_texture_idx[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_texture_idx[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_texture_idx")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetGlyphTextureIdx {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_glyph_texture_idx[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_glyph_texture_idx[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_glyph_texture_idx")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphTextureRid {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_texture_rid[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_texture_rid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_texture_rid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphTextureSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_texture_size[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_texture_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_texture_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphContours {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_contours[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_contours[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_contours")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetKerningList {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_kerning_list[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_kerning_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_kerning_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontClearKerningMap {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_clear_kerning_map[T](nil, nil, nil) } }

		func := textserverextension_gd_font_clear_kerning_map[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_clear_kerning_map")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRemoveKerning {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_remove_kerning[T](nil, nil, nil) } }

		func := textserverextension_gd_font_remove_kerning[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_remove_kerning")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetKerning {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_kerning[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_kerning[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_kerning")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetKerning {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_kerning[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_kerning[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_kerning")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlyphIndex {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_glyph_index[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_glyph_index[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_glyph_index")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetCharFromGlyphIndex {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_char_from_glyph_index[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_char_from_glyph_index[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_char_from_glyph_index")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontHasChar {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_has_char[T](nil, nil, nil) } }

		func := textserverextension_gd_font_has_char[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_has_char")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetSupportedChars {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_supported_chars[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_supported_chars[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_supported_chars")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetSupportedGlyphs {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_supported_glyphs[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_supported_glyphs[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_supported_glyphs")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRenderRange {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_render_range[T](nil, nil, nil) } }

		func := textserverextension_gd_font_render_range[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_render_range")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRenderGlyph {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_render_glyph[T](nil, nil, nil) } }

		func := textserverextension_gd_font_render_glyph[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_render_glyph")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontDrawGlyph {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_draw_glyph[T](nil, nil, nil) } }

		func := textserverextension_gd_font_draw_glyph[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_draw_glyph")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontDrawGlyphOutline {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_draw_glyph_outline[T](nil, nil, nil) } }

		func := textserverextension_gd_font_draw_glyph_outline[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_draw_glyph_outline")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontIsLanguageSupported {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_is_language_supported[T](nil, nil, nil) } }

		func := textserverextension_gd_font_is_language_supported[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_is_language_supported")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetLanguageSupportOverride {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_language_support_override[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_language_support_override[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_language_support_override")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetLanguageSupportOverride {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_language_support_override[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_language_support_override[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_language_support_override")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRemoveLanguageSupportOverride {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_remove_language_support_override[T](nil, nil, nil) } }

		func := textserverextension_gd_font_remove_language_support_override[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_remove_language_support_override")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetLanguageSupportOverrides {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_language_support_overrides[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_language_support_overrides[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_language_support_overrides")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontIsScriptSupported {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_is_script_supported[T](nil, nil, nil) } }

		func := textserverextension_gd_font_is_script_supported[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_is_script_supported")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetScriptSupportOverride {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_script_support_override[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_script_support_override[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_script_support_override")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetScriptSupportOverride {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_script_support_override[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_script_support_override[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_script_support_override")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontRemoveScriptSupportOverride {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_remove_script_support_override[T](nil, nil, nil) } }

		func := textserverextension_gd_font_remove_script_support_override[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_remove_script_support_override")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetScriptSupportOverrides {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_script_support_overrides[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_script_support_overrides[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_script_support_overrides")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetOpentypeFeatureOverrides {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_opentype_feature_overrides[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_opentype_feature_overrides[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_opentype_feature_overrides")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetOpentypeFeatureOverrides {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_opentype_feature_overrides[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_opentype_feature_overrides[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_opentype_feature_overrides")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSupportedFeatureList {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_supported_feature_list[T](nil, nil, nil) } }

		func := textserverextension_gd_font_supported_feature_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_supported_feature_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSupportedVariationList {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_supported_variation_list[T](nil, nil, nil) } }

		func := textserverextension_gd_font_supported_variation_list[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_supported_variation_list")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontGetGlobalOversampling {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_get_global_oversampling[T](nil, nil, nil) } }

		func := textserverextension_gd_font_get_global_oversampling[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_get_global_oversampling")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFontSetGlobalOversampling {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_font_set_global_oversampling[T](nil, nil, nil) } }

		func := textserverextension_gd_font_set_global_oversampling[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_font_set_global_oversampling")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionGetHexCodeBoxSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_get_hex_code_box_size[T](nil, nil, nil) } }

		func := textserverextension_gd_get_hex_code_box_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_hex_code_box_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionDrawHexCodeBox {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_draw_hex_code_box[T](nil, nil, nil) } }

		func := textserverextension_gd_draw_hex_code_box[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw_hex_code_box")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionCreateShapedText {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_create_shaped_text[T](nil, nil, nil) } }

		func := textserverextension_gd_create_shaped_text[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_shaped_text")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextClear {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_clear[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_clear[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_clear")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetDirection {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_direction[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_direction[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_direction")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetDirection {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_direction[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_direction[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_direction")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetInferredDirection {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_inferred_direction[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_inferred_direction[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_inferred_direction")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetBidiOverride {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_bidi_override[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_bidi_override[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_bidi_override")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetCustomPunctuation {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_custom_punctuation[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_custom_punctuation[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_custom_punctuation")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetCustomPunctuation {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_custom_punctuation[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_custom_punctuation[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_custom_punctuation")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetCustomEllipsis {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_custom_ellipsis[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_custom_ellipsis[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_custom_ellipsis")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetCustomEllipsis {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_custom_ellipsis[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_custom_ellipsis[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_custom_ellipsis")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetOrientation {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_orientation[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_orientation[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_orientation")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetOrientation {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_orientation[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_orientation[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_orientation")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetPreserveInvalid {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_preserve_invalid[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_preserve_invalid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_preserve_invalid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetPreserveInvalid {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_preserve_invalid[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_preserve_invalid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_preserve_invalid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetPreserveControl {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_preserve_control[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_preserve_control[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_preserve_control")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetPreserveControl {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_preserve_control[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_preserve_control[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_preserve_control")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSetSpacing {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_set_spacing[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_set_spacing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_set_spacing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetSpacing {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_spacing[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_spacing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_spacing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextAddString {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_add_string[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_add_string[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_add_string")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextAddObject {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_add_object[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_add_object[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_add_object")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextResizeObject {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_resize_object[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_resize_object[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_resize_object")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetText {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_text[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_text[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_text")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetSpanCount {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_span_count[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_span_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_span_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetSpanMeta {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_span_meta[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_span_meta[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_span_meta")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetSpanEmbeddedObject {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_span_embedded_object[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_span_embedded_object[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_span_embedded_object")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetSpanText {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_span_text[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_span_text[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_span_text")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetSpanObject {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_span_object[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_span_object[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_span_object")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedSetSpanUpdateFont {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_set_span_update_font[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_set_span_update_font[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_set_span_update_font")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunCount {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_count[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunText {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_text[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_text[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_text")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunRange {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_range[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_range[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_range")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunFontRid {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_font_rid[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_font_rid[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_font_rid")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunFontSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_font_size[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_font_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_font_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunLanguage {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_language[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_language[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_language")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunDirection {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_direction[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_direction[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_direction")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedGetRunObject {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_get_run_object[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_get_run_object[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_get_run_object")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSubstr {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_substr[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_substr[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_substr")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetParent {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_parent[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_parent[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_parent")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextFitToWidth {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_fit_to_width[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_fit_to_width[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_fit_to_width")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextTabAlign {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_tab_align[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_tab_align[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_tab_align")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextShape {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_shape[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_shape[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_shape")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextUpdateBreaks {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_update_breaks[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_update_breaks[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_update_breaks")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextUpdateJustificationOps {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_update_justification_ops[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_update_justification_ops[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_update_justification_ops")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextIsReady {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_is_ready[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_is_ready[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_is_ready")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetGlyphs {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_glyphs[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_glyphs[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_glyphs")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextSortLogical {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_sort_logical[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_sort_logical[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_sort_logical")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetGlyphCount {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_glyph_count[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_glyph_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_glyph_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetRange {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_range[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_range[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_range")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetLineBreaksAdv {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_line_breaks_adv[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_line_breaks_adv[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_line_breaks_adv")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetLineBreaks {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_line_breaks[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_line_breaks[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_line_breaks")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetWordBreaks {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_word_breaks[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_word_breaks[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_word_breaks")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetTrimPos {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_trim_pos[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_trim_pos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_trim_pos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetEllipsisPos {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_ellipsis_pos[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_ellipsis_pos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_ellipsis_pos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetEllipsisGlyphCount {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_ellipsis_glyph_count[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_ellipsis_glyph_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_ellipsis_glyph_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetEllipsisGlyphs {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_ellipsis_glyphs[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_ellipsis_glyphs[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_ellipsis_glyphs")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextOverrunTrimToWidth {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_overrun_trim_to_width[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_overrun_trim_to_width[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_overrun_trim_to_width")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetObjects {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_objects[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_objects[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_objects")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetObjectRect {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_object_rect[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_object_rect[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_object_rect")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetObjectRange {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_object_range[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_object_range[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_object_range")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetObjectGlyph {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_object_glyph[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_object_glyph[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_object_glyph")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetSize {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_size[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetAscent {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_ascent[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_ascent[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_ascent")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetDescent {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_descent[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_descent[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_descent")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetWidth {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_width[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_width[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_width")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetUnderlinePosition {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_underline_position[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_underline_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_underline_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetUnderlineThickness {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_underline_thickness[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_underline_thickness[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_underline_thickness")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetDominantDirectionInRange {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_dominant_direction_in_range[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_dominant_direction_in_range[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_dominant_direction_in_range")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetCarets {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_carets[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_carets[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_carets")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetSelection {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_selection[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_selection[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_selection")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextHitTestGrapheme {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_hit_test_grapheme[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_hit_test_grapheme[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_hit_test_grapheme")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextHitTestPosition {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_hit_test_position[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_hit_test_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_hit_test_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextDraw {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_draw[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_draw[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_draw")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextDrawOutline {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_draw_outline[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_draw_outline[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_draw_outline")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetGraphemeBounds {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_grapheme_bounds[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_grapheme_bounds[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_grapheme_bounds")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextNextGraphemePos {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_next_grapheme_pos[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_next_grapheme_pos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_next_grapheme_pos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextPrevGraphemePos {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_prev_grapheme_pos[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_prev_grapheme_pos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_prev_grapheme_pos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextGetCharacterBreaks {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_get_character_breaks[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_get_character_breaks[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_get_character_breaks")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextNextCharacterPos {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_next_character_pos[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_next_character_pos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_next_character_pos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextPrevCharacterPos {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_prev_character_pos[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_prev_character_pos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_prev_character_pos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionShapedTextClosestCharacterPos {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_shaped_text_closest_character_pos[T](nil, nil, nil) } }

		func := textserverextension_gd_shaped_text_closest_character_pos[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_shaped_text_closest_character_pos")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionFormatNumber {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_format_number[T](nil, nil, nil) } }

		func := textserverextension_gd_format_number[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_format_number")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionParseNumber {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_parse_number[T](nil, nil, nil) } }

		func := textserverextension_gd_parse_number[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_number")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionPercentSign {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_percent_sign[T](nil, nil, nil) } }

		func := textserverextension_gd_percent_sign[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_percent_sign")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionStripDiacritics {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_strip_diacritics[T](nil, nil, nil) } }

		func := textserverextension_gd_strip_diacritics[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_strip_diacritics")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionIsValidIdentifier {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_is_valid_identifier[T](nil, nil, nil) } }

		func := textserverextension_gd_is_valid_identifier[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_valid_identifier")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionIsValidLetter {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_is_valid_letter[T](nil, nil, nil) } }

		func := textserverextension_gd_is_valid_letter[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_valid_letter")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionStringGetWordBreaks {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_string_get_word_breaks[T](nil, nil, nil) } }

		func := textserverextension_gd_string_get_word_breaks[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_string_get_word_breaks")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionStringGetCharacterBreaks {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_string_get_character_breaks[T](nil, nil, nil) } }

		func := textserverextension_gd_string_get_character_breaks[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_string_get_character_breaks")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionIsConfusable {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_is_confusable[T](nil, nil, nil) } }

		func := textserverextension_gd_is_confusable[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_confusable")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionSpoofCheck {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_spoof_check[T](nil, nil, nil) } }

		func := textserverextension_gd_spoof_check[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_spoof_check")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionStringToUpper {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_string_to_upper[T](nil, nil, nil) } }

		func := textserverextension_gd_string_to_upper[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_string_to_upper")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionStringToLower {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_string_to_lower[T](nil, nil, nil) } }

		func := textserverextension_gd_string_to_lower[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_string_to_lower")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionStringToTitle {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_string_to_title[T](nil, nil, nil) } }

		func := textserverextension_gd_string_to_title[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_string_to_title")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionParseStructuredText {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_parse_structured_text[T](nil, nil, nil) } }

		func := textserverextension_gd_parse_structured_text[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_parse_structured_text")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextServerExtensionCleanup {{
		// HACK: force function generation
		if false { unsafe { textserverextension_gd_cleanup[T](nil, nil, nil) } }

		func := textserverextension_gd_cleanup[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_cleanup")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture2DGetWidth {{
		// HACK: force function generation
		if false { unsafe { texture2d_gd_get_width[T](nil, nil, nil) } }

		func := texture2d_gd_get_width[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_width")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture2DGetHeight {{
		// HACK: force function generation
		if false { unsafe { texture2d_gd_get_height[T](nil, nil, nil) } }

		func := texture2d_gd_get_height[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_height")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture2DIsPixelOpaque {{
		// HACK: force function generation
		if false { unsafe { texture2d_gd_is_pixel_opaque[T](nil, nil, nil) } }

		func := texture2d_gd_is_pixel_opaque[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_pixel_opaque")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture2DHasAlpha {{
		// HACK: force function generation
		if false { unsafe { texture2d_gd_has_alpha[T](nil, nil, nil) } }

		func := texture2d_gd_has_alpha[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_alpha")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture2DDraw {{
		// HACK: force function generation
		if false { unsafe { texture2d_gd_draw[T](nil, nil, nil) } }

		func := texture2d_gd_draw[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture2DDrawRect {{
		// HACK: force function generation
		if false { unsafe { texture2d_gd_draw_rect[T](nil, nil, nil) } }

		func := texture2d_gd_draw_rect[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw_rect")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture2DDrawRectRegion {{
		// HACK: force function generation
		if false { unsafe { texture2d_gd_draw_rect_region[T](nil, nil, nil) } }

		func := texture2d_gd_draw_rect_region[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_draw_rect_region")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture3DGetFormat {{
		// HACK: force function generation
		if false { unsafe { texture3d_gd_get_format[T](nil, nil, nil) } }

		func := texture3d_gd_get_format[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_format")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture3DGetWidth {{
		// HACK: force function generation
		if false { unsafe { texture3d_gd_get_width[T](nil, nil, nil) } }

		func := texture3d_gd_get_width[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_width")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture3DGetHeight {{
		// HACK: force function generation
		if false { unsafe { texture3d_gd_get_height[T](nil, nil, nil) } }

		func := texture3d_gd_get_height[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_height")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture3DGetDepth {{
		// HACK: force function generation
		if false { unsafe { texture3d_gd_get_depth[T](nil, nil, nil) } }

		func := texture3d_gd_get_depth[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_depth")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture3DHasMipmaps {{
		// HACK: force function generation
		if false { unsafe { texture3d_gd_has_mipmaps[T](nil, nil, nil) } }

		func := texture3d_gd_has_mipmaps[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_mipmaps")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITexture3DGetData {{
		// HACK: force function generation
		if false { unsafe { texture3d_gd_get_data[T](nil, nil, nil) } }

		func := texture3d_gd_get_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextureLayeredGetFormat {{
		// HACK: force function generation
		if false { unsafe { texturelayered_gd_get_format[T](nil, nil, nil) } }

		func := texturelayered_gd_get_format[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_format")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextureLayeredGetLayeredType {{
		// HACK: force function generation
		if false { unsafe { texturelayered_gd_get_layered_type[T](nil, nil, nil) } }

		func := texturelayered_gd_get_layered_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_layered_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextureLayeredGetWidth {{
		// HACK: force function generation
		if false { unsafe { texturelayered_gd_get_width[T](nil, nil, nil) } }

		func := texturelayered_gd_get_width[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_width")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextureLayeredGetHeight {{
		// HACK: force function generation
		if false { unsafe { texturelayered_gd_get_height[T](nil, nil, nil) } }

		func := texturelayered_gd_get_height[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_height")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextureLayeredGetLayers {{
		// HACK: force function generation
		if false { unsafe { texturelayered_gd_get_layers[T](nil, nil, nil) } }

		func := texturelayered_gd_get_layers[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_layers")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextureLayeredHasMipmaps {{
		// HACK: force function generation
		if false { unsafe { texturelayered_gd_has_mipmaps[T](nil, nil, nil) } }

		func := texturelayered_gd_has_mipmaps[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_has_mipmaps")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITextureLayeredGetLayerData {{
		// HACK: force function generation
		if false { unsafe { texturelayered_gd_get_layer_data[T](nil, nil, nil) } }

		func := texturelayered_gd_get_layer_data[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_layer_data")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITileMapUseTileDataRuntimeUpdate {{
		// HACK: force function generation
		if false { unsafe { tilemap_gd_use_tile_data_runtime_update[T](nil, nil, nil) } }

		func := tilemap_gd_use_tile_data_runtime_update[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_use_tile_data_runtime_update")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITileMapTileDataRuntimeUpdate {{
		// HACK: force function generation
		if false { unsafe { tilemap_gd_tile_data_runtime_update[T](nil, nil, nil) } }

		func := tilemap_gd_tile_data_runtime_update[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_tile_data_runtime_update")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITileMapLayerUseTileDataRuntimeUpdate {{
		// HACK: force function generation
		if false { unsafe { tilemaplayer_gd_use_tile_data_runtime_update[T](nil, nil, nil) } }

		func := tilemaplayer_gd_use_tile_data_runtime_update[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_use_tile_data_runtime_update")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITileMapLayerTileDataRuntimeUpdate {{
		// HACK: force function generation
		if false { unsafe { tilemaplayer_gd_tile_data_runtime_update[T](nil, nil, nil) } }

		func := tilemaplayer_gd_tile_data_runtime_update[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_tile_data_runtime_update")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITileMapLayerUpdateCells {{
		// HACK: force function generation
		if false { unsafe { tilemaplayer_gd_update_cells[T](nil, nil, nil) } }

		func := tilemaplayer_gd_update_cells[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_update_cells")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITranslationGetPluralMessage {{
		// HACK: force function generation
		if false { unsafe { translation_gd_get_plural_message[T](nil, nil, nil) } }

		func := translation_gd_get_plural_message[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_plural_message")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is ITranslationGetMessage {{
		// HACK: force function generation
		if false { unsafe { translation_gd_get_message[T](nil, nil, nil) } }

		func := translation_gd_get_message[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_message")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamInstantiatePlayback {{
		// HACK: force function generation
		if false { unsafe { videostream_gd_instantiate_playback[T](nil, nil, nil) } }

		func := videostream_gd_instantiate_playback[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_instantiate_playback")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackStop {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_stop[T](nil, nil, nil) } }

		func := videostreamplayback_gd_stop[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_stop")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackPlay {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_play[T](nil, nil, nil) } }

		func := videostreamplayback_gd_play[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_play")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackIsPlaying {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_is_playing[T](nil, nil, nil) } }

		func := videostreamplayback_gd_is_playing[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_playing")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackSetPaused {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_set_paused[T](nil, nil, nil) } }

		func := videostreamplayback_gd_set_paused[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_paused")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackIsPaused {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_is_paused[T](nil, nil, nil) } }

		func := videostreamplayback_gd_is_paused[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_paused")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackGetLength {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_get_length[T](nil, nil, nil) } }

		func := videostreamplayback_gd_get_length[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_length")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackGetPlaybackPosition {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_get_playback_position[T](nil, nil, nil) } }

		func := videostreamplayback_gd_get_playback_position[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_playback_position")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackSeek {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_seek[T](nil, nil, nil) } }

		func := videostreamplayback_gd_seek[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_seek")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackSetAudioTrack {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_set_audio_track[T](nil, nil, nil) } }

		func := videostreamplayback_gd_set_audio_track[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_audio_track")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackGetTexture {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_get_texture[T](nil, nil, nil) } }

		func := videostreamplayback_gd_get_texture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_texture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackUpdate {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_update[T](nil, nil, nil) } }

		func := videostreamplayback_gd_update[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_update")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackGetChannels {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_get_channels[T](nil, nil, nil) } }

		func := videostreamplayback_gd_get_channels[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_channels")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVideoStreamPlaybackGetMixRate {{
		// HACK: force function generation
		if false { unsafe { videostreamplayback_gd_get_mix_rate[T](nil, nil, nil) } }

		func := videostreamplayback_gd_get_mix_rate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_mix_rate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualInstance3DGetAabb {{
		// HACK: force function generation
		if false { unsafe { visualinstance3d_gd_get_aabb[T](nil, nil, nil) } }

		func := visualinstance3d_gd_get_aabb[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_aabb")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetName {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_name[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetDescription {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_description[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_description[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_description")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetCategory {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_category[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_category[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_category")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetReturnIconType {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_return_icon_type[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_return_icon_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_return_icon_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetInputPortCount {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_input_port_count[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_input_port_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_input_port_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetInputPortType {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_input_port_type[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_input_port_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_input_port_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetInputPortName {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_input_port_name[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_input_port_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_input_port_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetInputPortDefaultValue {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_input_port_default_value[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_input_port_default_value[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_input_port_default_value")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetDefaultInputPort {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_default_input_port[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_default_input_port[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_default_input_port")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetOutputPortCount {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_output_port_count[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_output_port_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_output_port_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetOutputPortType {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_output_port_type[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_output_port_type[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_output_port_type")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetOutputPortName {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_output_port_name[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_output_port_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_output_port_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetPropertyCount {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_property_count[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_property_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_property_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetPropertyName {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_property_name[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_property_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_property_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetPropertyDefaultIndex {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_property_default_index[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_property_default_index[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_property_default_index")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetPropertyOptions {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_property_options[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_property_options[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_property_options")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetCode {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_code[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetFuncCode {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_func_code[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_func_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_func_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomGetGlobalCode {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_get_global_code[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_get_global_code[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_global_code")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomIsHighend {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_is_highend[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_is_highend[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_highend")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IVisualShaderNodeCustomIsAvailable {{
		// HACK: force function generation
		if false { unsafe { visualshadernodecustom_gd_is_available[T](nil, nil, nil) } }

		func := visualshadernodecustom_gd_is_available[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_available")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetPacket {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_packet[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_packet[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_packet")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionPutPacket {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_put_packet[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_put_packet[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_put_packet")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetAvailablePacketCount {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_available_packet_count[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_available_packet_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_available_packet_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetMaxPacketSize {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_max_packet_size[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_max_packet_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_max_packet_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionPoll {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_poll[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_poll[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_poll")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionClose {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_close[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_close[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_close")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionSetWriteMode {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_set_write_mode[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_set_write_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_write_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetWriteMode {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_write_mode[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_write_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_write_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionWasStringPacket {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_was_string_packet[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_was_string_packet[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_was_string_packet")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetReadyState {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_ready_state[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_ready_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_ready_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetLabel {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_label[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_label[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_label")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionIsOrdered {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_is_ordered[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_is_ordered[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_ordered")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetId {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_id[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetMaxPacketLifeTime {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_max_packet_life_time[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_max_packet_life_time[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_max_packet_life_time")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetMaxRetransmits {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_max_retransmits[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_max_retransmits[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_max_retransmits")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetProtocol {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_protocol[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_protocol[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_protocol")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionIsNegotiated {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_is_negotiated[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_is_negotiated[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_negotiated")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCDataChannelExtensionGetBufferedAmount {{
		// HACK: force function generation
		if false { unsafe { webrtcdatachannelextension_gd_get_buffered_amount[T](nil, nil, nil) } }

		func := webrtcdatachannelextension_gd_get_buffered_amount[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_buffered_amount")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionGetConnectionState {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_get_connection_state[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_get_connection_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_connection_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionGetGatheringState {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_get_gathering_state[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_get_gathering_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_gathering_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionGetSignalingState {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_get_signaling_state[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_get_signaling_state[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_signaling_state")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionInitialize {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_initialize[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_initialize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_initialize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionCreateDataChannel {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_create_data_channel[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_create_data_channel[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_data_channel")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionCreateOffer {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_create_offer[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_create_offer[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_create_offer")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionSetRemoteDescription {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_set_remote_description[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_set_remote_description[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_remote_description")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionSetLocalDescription {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_set_local_description[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_set_local_description[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_local_description")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionAddIceCandidate {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_add_ice_candidate[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_add_ice_candidate[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_add_ice_candidate")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionPoll {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_poll[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_poll[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_poll")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWebRTCPeerConnectionExtensionClose {{
		// HACK: force function generation
		if false { unsafe { webrtcpeerconnectionextension_gd_close[T](nil, nil, nil) } }

		func := webrtcpeerconnectionextension_gd_close[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_close")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IWindowGetContentsMinimumSize {{
		// HACK: force function generation
		if false { unsafe { window_gd_get_contents_minimum_size[T](nil, nil, nil) } }

		func := window_gd_get_contents_minimum_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_contents_minimum_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetName {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_name[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_name[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_name")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetCapabilities {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_capabilities[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_capabilities[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_capabilities")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionIsInitialized {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_is_initialized[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_is_initialized[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_is_initialized")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionInitialize {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_initialize[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_initialize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_initialize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionUninitialize {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_uninitialize[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_uninitialize[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_uninitialize")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetSystemInfo {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_system_info[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_system_info[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_system_info")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionSupportsPlayAreaMode {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_supports_play_area_mode[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_supports_play_area_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_supports_play_area_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetPlayAreaMode {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_play_area_mode[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_play_area_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_play_area_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionSetPlayAreaMode {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_set_play_area_mode[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_set_play_area_mode[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_play_area_mode")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetPlayArea {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_play_area[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_play_area[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_play_area")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetRenderTargetSize {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_render_target_size[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_render_target_size[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_render_target_size")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetViewCount {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_view_count[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_view_count[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_view_count")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetCameraTransform {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_camera_transform[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_camera_transform[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_camera_transform")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetTransformForView {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_transform_for_view[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_transform_for_view[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_transform_for_view")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetProjectionForView {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_projection_for_view[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_projection_for_view[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_projection_for_view")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetVrsTexture {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_vrs_texture[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_vrs_texture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_vrs_texture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionProcess {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_process[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_process[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_process")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionPreRender {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_pre_render[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_pre_render[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pre_render")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionPreDrawViewport {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_pre_draw_viewport[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_pre_draw_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_pre_draw_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionPostDrawViewport {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_post_draw_viewport[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_post_draw_viewport[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_post_draw_viewport")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionEndFrame {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_end_frame[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_end_frame[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_end_frame")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetSuggestedTrackerNames {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_suggested_tracker_names[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_suggested_tracker_names[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_suggested_tracker_names")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetSuggestedPoseNames {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_suggested_pose_names[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_suggested_pose_names[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_suggested_pose_names")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetTrackingStatus {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_tracking_status[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_tracking_status[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_tracking_status")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionTriggerHapticPulse {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_trigger_haptic_pulse[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_trigger_haptic_pulse[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_trigger_haptic_pulse")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetAnchorDetectionIsEnabled {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_anchor_detection_is_enabled[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_anchor_detection_is_enabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_anchor_detection_is_enabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionSetAnchorDetectionIsEnabled {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_set_anchor_detection_is_enabled[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_set_anchor_detection_is_enabled[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_set_anchor_detection_is_enabled")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetCameraFeedId {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_camera_feed_id[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_camera_feed_id[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_camera_feed_id")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetColorTexture {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_color_texture[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_color_texture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_color_texture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetDepthTexture {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_depth_texture[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_depth_texture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_depth_texture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
	$if T is IXRInterfaceExtensionGetVelocityTexture {{
		// HACK: force function generation
		if false { unsafe { xrinterfaceextension_gd_get_velocity_texture[T](nil, nil, nil) } }

		func := xrinterfaceextension_gd_get_velocity_texture[T]
		ivar := i64(func)
		var := i64_to_variant(ivar)
		sn := StringName.new("_get_velocity_texture")
		ci.virtual_methods.index_set_named(sn, var) or {panic(err)}
		sn.deinit()
	}}
}
