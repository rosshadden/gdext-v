module gd

pub struct MenuButton {
	Button
}

pub fn (s &MenuButton) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s MenuButton) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &MenuButton) get_popup() PopupMenu {
	mut result := PopupMenu{}
	classname := StringName.new("MenuButton")
	fnname := StringName.new("get_popup")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 229722558)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &MenuButton) show_popup() {
	classname := StringName.new("MenuButton")
	fnname := StringName.new("show_popup")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &MenuButton) set_switch_on_hover(enable bool) {
	classname := StringName.new("MenuButton")
	fnname := StringName.new("set_switch_on_hover")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&enable)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &MenuButton) is_switch_on_hover() bool {
	mut result := false
	classname := StringName.new("MenuButton")
	fnname := StringName.new("is_switch_on_hover")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2240911060)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &MenuButton) set_disable_shortcuts(disabled bool) {
	classname := StringName.new("MenuButton")
	fnname := StringName.new("set_disable_shortcuts")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&disabled)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &MenuButton) set_item_count(count i64) {
	classname := StringName.new("MenuButton")
	fnname := StringName.new("set_item_count")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&count)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &MenuButton) get_item_count() i64 {
	mut result := i64(0)
	classname := StringName.new("MenuButton")
	fnname := StringName.new("get_item_count")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
