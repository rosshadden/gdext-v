module gd

pub struct AnimationNodeTimeSeek {
	AnimationNode
}

pub fn (s &AnimationNodeTimeSeek) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s AnimationNodeTimeSeek) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &AnimationNodeTimeSeek) set_explicit_elapse(enable bool) {
	classname := StringName.new("AnimationNodeTimeSeek")
	fnname := StringName.new("set_explicit_elapse")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&enable)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &AnimationNodeTimeSeek) is_explicit_elapse() bool {
	mut result := false
	classname := StringName.new("AnimationNodeTimeSeek")
	fnname := StringName.new("is_explicit_elapse")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
