module gd

pub struct ParallaxLayer {
	Node2D
}

pub fn (s &ParallaxLayer) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s ParallaxLayer) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &ParallaxLayer) set_motion_scale(scale Vector2) {
	classname := StringName.new("ParallaxLayer")
	fnname := StringName.new("set_motion_scale")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 743155724)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&scale)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &ParallaxLayer) get_motion_scale() Vector2 {
	mut result := Vector2{}
	classname := StringName.new("ParallaxLayer")
	fnname := StringName.new("get_motion_scale")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &ParallaxLayer) set_motion_offset(offset Vector2) {
	classname := StringName.new("ParallaxLayer")
	fnname := StringName.new("set_motion_offset")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 743155724)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&offset)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &ParallaxLayer) get_motion_offset() Vector2 {
	mut result := Vector2{}
	classname := StringName.new("ParallaxLayer")
	fnname := StringName.new("get_motion_offset")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &ParallaxLayer) set_mirroring(mirror Vector2) {
	classname := StringName.new("ParallaxLayer")
	fnname := StringName.new("set_mirroring")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 743155724)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&mirror)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &ParallaxLayer) get_mirroring() Vector2 {
	mut result := Vector2{}
	classname := StringName.new("ParallaxLayer")
	fnname := StringName.new("get_mirroring")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
