module gd

pub struct MultiMeshInstance3D {
	GeometryInstance3D
}

pub fn (s &MultiMeshInstance3D) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s MultiMeshInstance3D) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &MultiMeshInstance3D) set_multimesh(multimesh MultiMesh) {
	classname := StringName.new("MultiMeshInstance3D")
	fnname := StringName.new("set_multimesh")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2246127404)
	mut args := unsafe { [1]voidptr{} }
	args[0] = voidptr(&multimesh.ptr)
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &MultiMeshInstance3D) get_multimesh() MultiMesh {
	mut result := MultiMesh{}
	classname := StringName.new("MultiMeshInstance3D")
	fnname := StringName.new("get_multimesh")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1385450523)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}
