module gd

pub struct TranslationServer {
	Object
}

pub fn TranslationServer.get_singleton() TranslationServer {
	sn := StringName.new("TranslationServer")
	result := TranslationServer{
		ptr: gdf.global_get_singleton(sn)
	}
	sn.deinit()
	return result
}

pub fn (s &TranslationServer) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s TranslationServer) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

pub fn (s &TranslationServer) set_locale(locale string) {
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("set_locale")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 83702148)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := String.new(locale)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
}

pub fn (s &TranslationServer) get_locale() string {
	mut result := String{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_locale")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 201670096)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &TranslationServer) get_tool_locale() string {
	mut result := String{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_tool_locale")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2841200299)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &TranslationServer) compare_locales(locale_a string, locale_b string) i64 {
	mut result := i64(0)
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("compare_locales")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2878152881)
	mut args := unsafe { [2]voidptr{} }
	arg_sn0 := String.new(locale_a)
	args[0] = unsafe{voidptr(&arg_sn0)}
	arg_sn1 := String.new(locale_b)
	args[1] = unsafe{voidptr(&arg_sn1)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	arg_sn1.deinit()
	classname.deinit()
	fnname.deinit()
	return result
}

@[params]
pub struct TranslationServer_standardize_locale_Cfg {
pub:
	add_defaults bool
}

pub fn (s &TranslationServer) standardize_locale(locale string, cfg TranslationServer_standardize_locale_Cfg) string {
	mut result := String{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("standardize_locale")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 4216441673)
	mut args := unsafe { [2]voidptr{} }
	arg_sn0 := String.new(locale)
	args[0] = unsafe{voidptr(&arg_sn0)}
	args[1] = unsafe{voidptr(&cfg.add_defaults)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &TranslationServer) get_all_languages() PackedStringArray {
	mut result := PackedStringArray{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_all_languages")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1139954409)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) get_language_name(language string) string {
	mut result := String{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_language_name")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3135753539)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := String.new(language)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &TranslationServer) get_all_scripts() PackedStringArray {
	mut result := PackedStringArray{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_all_scripts")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1139954409)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) get_script_name(script string) string {
	mut result := String{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_script_name")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3135753539)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := String.new(script)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &TranslationServer) get_all_countries() PackedStringArray {
	mut result := PackedStringArray{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_all_countries")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1139954409)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) get_country_name(country string) string {
	mut result := String{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_country_name")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3135753539)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := String.new(country)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &TranslationServer) get_locale_name(locale string) string {
	mut result := String{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_locale_name")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3135753539)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := String.new(locale)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

@[params]
pub struct TranslationServer_translate_Cfg {
pub:
	context string
}

pub fn (s &TranslationServer) translate(message string, cfg TranslationServer_translate_Cfg) string {
	mut result := StringName{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("translate")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1829228469)
	mut args := unsafe { [2]voidptr{} }
	arg_sn0 := StringName.new(message)
	args[0] = unsafe{voidptr(&arg_sn0)}
	arg_sn1 := StringName.new(cfg.context)
	args[1] = unsafe{voidptr(&arg_sn1)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	arg_sn1.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

@[params]
pub struct TranslationServer_translate_plural_Cfg {
pub:
	context string
}

pub fn (s &TranslationServer) translate_plural(message string, plural_message string, n i64, cfg TranslationServer_translate_plural_Cfg) string {
	mut result := StringName{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("translate_plural")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 229954002)
	mut args := unsafe { [4]voidptr{} }
	arg_sn0 := StringName.new(message)
	args[0] = unsafe{voidptr(&arg_sn0)}
	arg_sn1 := StringName.new(plural_message)
	args[1] = unsafe{voidptr(&arg_sn1)}
	args[2] = unsafe{voidptr(&n)}
	arg_sn3 := StringName.new(cfg.context)
	args[3] = unsafe{voidptr(&arg_sn3)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	arg_sn1.deinit()
	arg_sn3.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &TranslationServer) add_translation(translation Translation) {
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("add_translation")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1466479800)
	mut args := unsafe { [1]voidptr{} }
	args[0] = voidptr(&translation.ptr)
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &TranslationServer) remove_translation(translation Translation) {
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("remove_translation")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1466479800)
	mut args := unsafe { [1]voidptr{} }
	args[0] = voidptr(&translation.ptr)
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &TranslationServer) get_translation_object(locale string) Translation {
	mut result := Translation{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_translation_object")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2065240175)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := String.new(locale)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) has_domain(domain string) bool {
	mut result := false
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("has_domain")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2619796661)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := StringName.new(domain)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) get_or_add_domain(domain string) TranslationDomain {
	mut result := TranslationDomain{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_or_add_domain")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 397200075)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := StringName.new(domain)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) remove_domain(domain string) {
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("remove_domain")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3304788590)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := StringName.new(domain)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
}

pub fn (s &TranslationServer) clear() {
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("clear")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &TranslationServer) get_loaded_locales() PackedStringArray {
	mut result := PackedStringArray{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("get_loaded_locales")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1139954409)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) is_pseudolocalization_enabled() bool {
	mut result := false
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("is_pseudolocalization_enabled")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &TranslationServer) set_pseudolocalization_enabled(enabled bool) {
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("set_pseudolocalization_enabled")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&enabled)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &TranslationServer) reload_pseudolocalization() {
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("reload_pseudolocalization")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &TranslationServer) pseudolocalize(message string) string {
	mut result := StringName{}
	classname := StringName.new("TranslationServer")
	fnname := StringName.new("pseudolocalize")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1965194235)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := StringName.new(message)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}
