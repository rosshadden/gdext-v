module gd

// TODO: this will be generated from the API dump in _GDExtension.v, once enums are mapped
pub enum GDExtensionInitializationLevel as i64 {
	initialization_level_core    = 0
	initialization_level_servers = 1
	initialization_level_scene   = 2
	initialization_level_editor  = 3
}
