module gd

pub struct OptionButton {
	Button
}

pub fn (s &OptionButton) to_variant() Variant {
	to_variant := gdf.get_variant_from_type_constructor(GDExtensionVariantType.type_object)
	result := Variant{}
	to_variant(GDExtensionUninitializedVariantPtr(&result), s.ptr)
	return result
}

pub fn (mut s OptionButton) from_variant(var &Variant) {
	variant_to_type := gdf.get_variant_to_type_constructor(GDExtensionVariantType.type_object)
	variant_to_type(voidptr(&s.ptr), var)
}

@[params]
pub struct OptionButton_add_item_Cfg {
pub:
	id i64
}

pub fn (s &OptionButton) add_item(label string, cfg OptionButton_add_item_Cfg) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("add_item")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2697778442)
	mut args := unsafe { [2]voidptr{} }
	arg_sn0 := String.new(label)
	args[0] = unsafe{voidptr(&arg_sn0)}
	args[1] = unsafe{voidptr(&cfg.id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
}

@[params]
pub struct OptionButton_add_icon_item_Cfg {
pub:
	id i64
}

pub fn (s &OptionButton) add_icon_item(texture Texture2D, label string, cfg OptionButton_add_icon_item_Cfg) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("add_icon_item")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3781678508)
	mut args := unsafe { [3]voidptr{} }
	args[0] = voidptr(&texture.ptr)
	arg_sn1 := String.new(label)
	args[1] = unsafe{voidptr(&arg_sn1)}
	args[2] = unsafe{voidptr(&cfg.id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn1.deinit()
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_text(idx i64, text string) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_text")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 501894301)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	arg_sn1 := String.new(text)
	args[1] = unsafe{voidptr(&arg_sn1)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn1.deinit()
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_icon(idx i64, texture Texture2D) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_icon")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 666127730)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	args[1] = voidptr(&texture.ptr)
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_disabled(idx i64, disabled bool) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_disabled")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 300928843)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	args[1] = unsafe{voidptr(&disabled)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_id(idx i64, id i64) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_id")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3937882851)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	args[1] = unsafe{voidptr(&id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_metadata(idx i64, metadata Variant) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_metadata")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2152698145)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	args[1] = unsafe{voidptr(&metadata)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_tooltip(idx i64, tooltip string) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_tooltip")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 501894301)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	arg_sn1 := String.new(tooltip)
	args[1] = unsafe{voidptr(&arg_sn1)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn1.deinit()
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_auto_translate_mode(idx i64, mode NodeAutoTranslateMode) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_auto_translate_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 287402019)
	mut args := unsafe { [2]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	i64_mode := i64(mode)
	args[1] = unsafe{voidptr(&i64_mode)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) get_item_text(idx i64) string {
	mut result := String{}
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_text")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 844755477)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &OptionButton) get_item_icon(idx i64) Texture2D {
	mut result := Texture2D{}
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_icon")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3536238170)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) get_item_id(idx i64) i64 {
	mut result := i64(0)
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_id")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 923996154)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) get_item_index(id i64) i64 {
	mut result := i64(0)
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_index")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 923996154)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&id)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) get_item_metadata(idx i64) Variant {
	mut result := Variant{}
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_metadata")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 4227898402)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) get_item_tooltip(idx i64) string {
	mut result := String{}
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_tooltip")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 844755477)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	result_v := result.to_v()
	result.deinit()
	return result_v
}

pub fn (s &OptionButton) get_item_auto_translate_mode(idx i64) NodeAutoTranslateMode {
	mut result := i64(NodeAutoTranslateMode.auto_translate_mode_inherit)
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_auto_translate_mode")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 906302372)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return unsafe{NodeAutoTranslateMode(result)}
}

pub fn (s &OptionButton) is_item_disabled(idx i64) bool {
	mut result := false
	classname := StringName.new("OptionButton")
	fnname := StringName.new("is_item_disabled")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1116898809)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) is_item_separator(idx i64) bool {
	mut result := false
	classname := StringName.new("OptionButton")
	fnname := StringName.new("is_item_separator")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1116898809)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

@[params]
pub struct OptionButton_add_separator_Cfg {
pub:
	text string
}

pub fn (s &OptionButton) add_separator(cfg OptionButton_add_separator_Cfg) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("add_separator")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3005725572)
	mut args := unsafe { [1]voidptr{} }
	arg_sn0 := String.new(cfg.text)
	args[0] = unsafe{voidptr(&arg_sn0)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	arg_sn0.deinit()
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) clear() {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("clear")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) gd_select(idx i64) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("select")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) get_selected() i64 {
	mut result := i64(0)
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_selected")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) get_selected_id() i64 {
	mut result := i64(0)
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_selected_id")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) get_selected_metadata() Variant {
	mut result := Variant{}
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_selected_metadata")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1214101251)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) remove_item(idx i64) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("remove_item")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&idx)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) get_popup() PopupMenu {
	mut result := PopupMenu{}
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_popup")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 229722558)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) show_popup() {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("show_popup")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) set_item_count(count i64) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_item_count")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 1286410249)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&count)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) get_item_count() i64 {
	mut result := i64(0)
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_item_count")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) has_selectable_items() bool {
	mut result := false
	classname := StringName.new("OptionButton")
	fnname := StringName.new("has_selectable_items")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

@[params]
pub struct OptionButton_get_selectable_item_Cfg {
pub:
	from_last bool
}

pub fn (s &OptionButton) get_selectable_item(cfg OptionButton_get_selectable_item_Cfg) i64 {
	mut result := i64(0)
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_selectable_item")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 894402480)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&cfg.from_last)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) set_fit_to_longest_item(fit bool) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_fit_to_longest_item")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&fit)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) is_fit_to_longest_item() bool {
	mut result := false
	classname := StringName.new("OptionButton")
	fnname := StringName.new("is_fit_to_longest_item")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) set_allow_reselect(allow bool) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_allow_reselect")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&allow)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}

pub fn (s &OptionButton) get_allow_reselect() bool {
	mut result := false
	classname := StringName.new("OptionButton")
	fnname := StringName.new("get_allow_reselect")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
	gdf.object_method_bind_ptrcall(mb, s.ptr, unsafe{nil}, voidptr(&result))
	classname.deinit()
	fnname.deinit()
	return result
}

pub fn (s &OptionButton) set_disable_shortcuts(disabled bool) {
	classname := StringName.new("OptionButton")
	fnname := StringName.new("set_disable_shortcuts")
	mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
	mut args := unsafe { [1]voidptr{} }
	args[0] = unsafe{voidptr(&disabled)}
	gdf.object_method_bind_ptrcall(mb, s.ptr, voidptr(&args[0]), unsafe{nil})
	classname.deinit()
	fnname.deinit()
}
